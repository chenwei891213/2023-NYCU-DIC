.title measure EDP
.vec 'Pattern_comparator.vec'
.include '../../16mos.pm'
.include '../../7nm_TT.pm'
.include '/RAID2/COURSE/dic/dic098/lab4/4-1/EDPMeasure/asap7sc7p5t_AO_RVT.sp'
.include '/RAID2/COURSE/dic/dic098/lab4/4-1/EDPMeasure/asap7sc7p5t_INVBUF_RVT.sp'
.include '/RAID2/COURSE/dic/dic098/lab4/4-1/EDPMeasure/asap7sc7p5t_OA_RVT.sp'
.include '/RAID2/COURSE/dic/dic098/lab4/4-1/EDPMeasure/asap7sc7p5t_SEQ_RVT.sp'
.include '/RAID2/COURSE/dic/dic098/lab4/4-1/EDPMeasure/asap7sc7p5t_SIMPLE_RVT.sp'
.include 'Comparator_SYN_new.sp'
* .include 'Original_Comparator_SYN_new.sp'
.param Vin = 0.4
VDD VDD GND  Vin
VSS VSS GND 0 

X1 VSS VDD  a0 a1 a2 a3 a4 a5 a6 a7 a8 a9  a10	a11	a12	a13	a14	a15	a16	a17	a18	a19	a20	a21	a22	a23	a24	a25	a26	a27	a28	a29	a30	a31	a32	a33	a34	a35	a36	a37	a38	a39	a40	a41	a42	a43	a44	a45	a46	a47	a48	a49	a50	a51	a52	a53	a54	a55	a56	a57	a58	a59	a60	a61	a62	a63 b0 b1 b2 b3 b4 b5 b6 b7 b8 b9	b10	b11	b12	b13	b14	b15	b16	b17	b18	b19	b20	b21	b22	b23	b24	b25	b26	b27	b28	b29	b30	b31	b32	b33	b34	b35	b36	b37	b38	b39	b40	b41	b42	b43	b44	b45	b46	b47	b48	b49	b50	b51	b52	b53	b54	b55	b56	b57	b58	b59	b60	b61	b62	b63 Out Comparator
X2 0 VDD a1 inv_a1 BUFX10_ASAP7_75T_R
X3 0 VDD a2 inv_a2 BUFX10_ASAP7_75T_R
X4 0 VDD a3 inv_a3 BUFX10_ASAP7_75T_R
X5 0 VDD a4 inv_a4 BUFX10_ASAP7_75T_R
X6 0 VDD a5 inv_a5 BUFX10_ASAP7_75T_R
X7 0 VDD a6 inv_a6 BUFX10_ASAP7_75T_R
X8 0 VDD a7 inv_a7 BUFX10_ASAP7_75T_R
X9 0 VDD a8 inv_a8 BUFX10_ASAP7_75T_R
X10 0 VDD a9 inv_a9 BUFX10_ASAP7_75T_R
X11 0 VDD a10 inv_a10 BUFX10_ASAP7_75T_R
X12 0 VDD a11 inv_a11 BUFX10_ASAP7_75T_R
X13 0 VDD a12 inv_a12 BUFX10_ASAP7_75T_R
X14 0 VDD a13 inv_a13 BUFX10_ASAP7_75T_R
X15 0 VDD a14 inv_a14 BUFX10_ASAP7_75T_R
X16 0 VDD a15 inv_a15 BUFX10_ASAP7_75T_R
X17 0 VDD a16 inv_a16 BUFX10_ASAP7_75T_R
X18 0 VDD a17 inv_a17 BUFX10_ASAP7_75T_R
X19 0 VDD a18 inv_a18 BUFX10_ASAP7_75T_R
X20 0 VDD a19 inv_a19 BUFX10_ASAP7_75T_R
X21 0 VDD a20 inv_a20 BUFX10_ASAP7_75T_R
X22 0 VDD a21 inv_a21 BUFX10_ASAP7_75T_R
X23 0 VDD a22 inv_a22 BUFX10_ASAP7_75T_R
X24 0 VDD a23 inv_a23 BUFX10_ASAP7_75T_R
X25 0 VDD a24 inv_a24 BUFX10_ASAP7_75T_R
X26 0 VDD a25 inv_a25 BUFX10_ASAP7_75T_R
X27 0 VDD a26 inv_a26 BUFX10_ASAP7_75T_R
X28 0 VDD a27 inv_a27 BUFX10_ASAP7_75T_R
X29 0 VDD a28 inv_a28 BUFX10_ASAP7_75T_R
X30 0 VDD a29 inv_a29 BUFX10_ASAP7_75T_R
X31 0 VDD a30 inv_a30 BUFX10_ASAP7_75T_R
X32 0 VDD a31 inv_a31 BUFX10_ASAP7_75T_R
X33 0 VDD a32 inv_a32 BUFX10_ASAP7_75T_R
X34 0 VDD a33 inv_a33 BUFX10_ASAP7_75T_R
X35 0 VDD a34 inv_a34 BUFX10_ASAP7_75T_R
X36 0 VDD a35 inv_a35 BUFX10_ASAP7_75T_R
X37 0 VDD a36 inv_a36 BUFX10_ASAP7_75T_R
X38 0 VDD a37 inv_a37 BUFX10_ASAP7_75T_R
X39 0 VDD a38 inv_a38 BUFX10_ASAP7_75T_R
X40 0 VDD a39 inv_a39 BUFX10_ASAP7_75T_R
X41 0 VDD a40 inv_a40 BUFX10_ASAP7_75T_R
X42 0 VDD a41 inv_a41 BUFX10_ASAP7_75T_R
X43 0 VDD a42 inv_a42 BUFX10_ASAP7_75T_R
X44 0 VDD a43 inv_a43 BUFX10_ASAP7_75T_R
X45 0 VDD a44 inv_a44 BUFX10_ASAP7_75T_R
X46 0 VDD a45 inv_a45 BUFX10_ASAP7_75T_R
X47 0 VDD a46 inv_a46 BUFX10_ASAP7_75T_R
X48 0 VDD a47 inv_a47 BUFX10_ASAP7_75T_R
X49 0 VDD a48 inv_a48 BUFX10_ASAP7_75T_R
X50 0 VDD a49 inv_a49 BUFX10_ASAP7_75T_R
X51 0 VDD a50 inv_a50 BUFX10_ASAP7_75T_R
X52 0 VDD a51 inv_a51 BUFX10_ASAP7_75T_R
X53 0 VDD a52 inv_a52 BUFX10_ASAP7_75T_R
X54 0 VDD a53 inv_a53 BUFX10_ASAP7_75T_R
X55 0 VDD a54 inv_a54 BUFX10_ASAP7_75T_R
X56 0 VDD a55 inv_a55 BUFX10_ASAP7_75T_R
X57 0 VDD a56 inv_a56 BUFX10_ASAP7_75T_R
X58 0 VDD a57 inv_a57 BUFX10_ASAP7_75T_R
X59 0 VDD a58 inv_a58 BUFX10_ASAP7_75T_R
X60 0 VDD a59 inv_a59 BUFX10_ASAP7_75T_R
X61 0 VDD a60 inv_a60 BUFX10_ASAP7_75T_R
X62 0 VDD a61 inv_a61 BUFX10_ASAP7_75T_R
X63 0 VDD a62 inv_a62 BUFX10_ASAP7_75T_R
X64 0 VDD b1 inv_b1 BUFX10_ASAP7_75T_R
X65 0 VDD b2 inv_b2 BUFX10_ASAP7_75T_R
X66 0 VDD b3 inv_b3 BUFX10_ASAP7_75T_R
X67 0 VDD b4 inv_b4 BUFX10_ASAP7_75T_R
X68 0 VDD b5 inv_b5 BUFX10_ASAP7_75T_R
X69 0 VDD b6 inv_b6 BUFX10_ASAP7_75T_R
X70 0 VDD b7 inv_b7 BUFX10_ASAP7_75T_R
X71 0 VDD b8 inv_b8 BUFX10_ASAP7_75T_R
X72 0 VDD b9 inv_b9 BUFX10_ASAP7_75T_R
X73 0 VDD b10 inv_b10 BUFX10_ASAP7_75T_R
X74 0 VDD b11 inv_b11 BUFX10_ASAP7_75T_R
X75 0 VDD b12 inv_b12 BUFX10_ASAP7_75T_R
X76 0 VDD b13 inv_b13 BUFX10_ASAP7_75T_R
X77 0 VDD b14 inv_b14 BUFX10_ASAP7_75T_R
X78 0 VDD b15 inv_b15 BUFX10_ASAP7_75T_R
X79 0 VDD b16 inv_b16 BUFX10_ASAP7_75T_R
X80 0 VDD b17 inv_b17 BUFX10_ASAP7_75T_R
X81 0 VDD b18 inv_b18 BUFX10_ASAP7_75T_R
X82 0 VDD b19 inv_b19 BUFX10_ASAP7_75T_R
X83 0 VDD b20 inv_b20 BUFX10_ASAP7_75T_R
X84 0 VDD b21 inv_b21 BUFX10_ASAP7_75T_R
X85 0 VDD b22 inv_b22 BUFX10_ASAP7_75T_R
X86 0 VDD b23 inv_b23 BUFX10_ASAP7_75T_R
X87 0 VDD b24 inv_b24 BUFX10_ASAP7_75T_R
X88 0 VDD b25 inv_b25 BUFX10_ASAP7_75T_R
X89 0 VDD b26 inv_b26 BUFX10_ASAP7_75T_R
X90 0 VDD b27 inv_b27 BUFX10_ASAP7_75T_R
X91 0 VDD b28 inv_b28 BUFX10_ASAP7_75T_R
X92 0 VDD b29 inv_b29 BUFX10_ASAP7_75T_R
X93 0 VDD b30 inv_b30 BUFX10_ASAP7_75T_R
X94 0 VDD b31 inv_b31 BUFX10_ASAP7_75T_R
X95 0 VDD b32 inv_b32 BUFX10_ASAP7_75T_R
X96 0 VDD b33 inv_b33 BUFX10_ASAP7_75T_R
X97 0 VDD b34 inv_b34 BUFX10_ASAP7_75T_R
X98 0 VDD b35 inv_b35 BUFX10_ASAP7_75T_R
X99 0 VDD b36 inv_b36 BUFX10_ASAP7_75T_R
X100 0 VDD b37 inv_b37 BUFX10_ASAP7_75T_R
X101 0 VDD b38 inv_b38 BUFX10_ASAP7_75T_R
X102 0 VDD b39 inv_b39 BUFX10_ASAP7_75T_R
X103 0 VDD b40 inv_b40 BUFX10_ASAP7_75T_R
X104 0 VDD b41 inv_b41 BUFX10_ASAP7_75T_R
X105 0 VDD b42 inv_b42 BUFX10_ASAP7_75T_R
X106 0 VDD b43 inv_b43 BUFX10_ASAP7_75T_R
X107 0 VDD b44 inv_b44 BUFX10_ASAP7_75T_R
X108 0 VDD b45 inv_b45 BUFX10_ASAP7_75T_R
X109 0 VDD b46 inv_b46 BUFX10_ASAP7_75T_R
X110 0 VDD b47 inv_b47 BUFX10_ASAP7_75T_R
X111 0 VDD b48 inv_b48 BUFX10_ASAP7_75T_R
X112 0 VDD b49 inv_b49 BUFX10_ASAP7_75T_R
X113 0 VDD b50 inv_b50 BUFX10_ASAP7_75T_R
X114 0 VDD b51 inv_b51 BUFX10_ASAP7_75T_R
X115 0 VDD b52 inv_b52 BUFX10_ASAP7_75T_R
X116 0 VDD b53 inv_b53 BUFX10_ASAP7_75T_R
X117 0 VDD b54 inv_b54 BUFX10_ASAP7_75T_R
X118 0 VDD b55 inv_b55 BUFX10_ASAP7_75T_R
X119 0 VDD b56 inv_b56 BUFX10_ASAP7_75T_R
X120 0 VDD b57 inv_b57 BUFX10_ASAP7_75T_R
X121 0 VDD b58 inv_b58 BUFX10_ASAP7_75T_R
X122 0 VDD b59 inv_b59 BUFX10_ASAP7_75T_R
X123 0 VDD b60 inv_b60 BUFX10_ASAP7_75T_R
X124 0 VDD b61 inv_b61 BUFX10_ASAP7_75T_R
X125 0 VDD b62 inv_b62 BUFX10_ASAP7_75T_R
X126 0 VDD a0 inv_a0 BUFX10_ASAP7_75T_R
X127 0 VDD a63 inv_a63 BUFX10_ASAP7_75T_R
X128 0 VDD b0 inv_b0 BUFX10_ASAP7_75T_R
X129 0 VDD b63 inv_b63 BUFX10_ASAP7_75T_R
Cout_loading out gnd 5fF
* Cwire_loading out gnd 3fF

* C2 Output[8] gnd 5fF
* C3 Output[7] gnd 5fF
* C4 Output[6] gnd 5fF
* C5 Output[5] gnd 5fF
* C6 Output[4] gnd 5fF
* C7 Output[3] gnd 5fF
* C8 Output[2] gnd 5fF
* C9 Output[1] gnd 5fF
* C0 Output[0] gnd 5fF
.tran 1ns 50*100ns 

.meas TRAN Delay TRIG V(a0) VAL=Vin/2 RISE=1
+TARG V(out) VAL = Vin/2 RISE=1
.meas TRAN Tr TRIG V(out) VAL=Vin*0.1 RISE=1
+TARG V(out) VAL = Vin*0.9 RISE=1
.meas TRAN Tf TRIG V(out) VAL=Vin*0.9 FALL=1
+TARG V(out) VAL = Vin*0.1 FALL=1
.measure TRAN Power avg  P(X1) from=0.0n to=50*100ns 
* .measure tran Energy INTEG V(VDD)*I(X1) FROM=0 TO=70us
.options post
.end
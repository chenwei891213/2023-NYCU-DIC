.SUBCKT Adder_4bit VSS VDD  A[3] A[2] A[1] A[0] B[3] B[2] B[1] B[0] Output[4] Output[3] Output[2] Output[1] Output[0]
XU3 VSS VDD  A[0] B[0] Output[0] XOR2xp5_ASAP7_75t_R
XU4 VSS VDD  B[0] A[0] n11 NAND2xp5_ASAP7_75t_R
XU5 VSS VDD  B[1] A[1] n11 A0  Output[1] FAx1_ASAP7_75t_R
XU6 VSS VDD  B[2] A[2] n6 XNOR2xp5_ASAP7_75t_R
XU7 VSS VDD  B[1] A[1] n9 NAND2xp5_ASAP7_75t_R
XU8 VSS VDD  n11 n9 n4 NAND2xp5_ASAP7_75t_R
XU9 VSS VDD  B[1] A[1] n7 OR2x2_ASAP7_75t_R
XU10 VSS VDD  n4 n7 n5 NAND2xp5_ASAP7_75t_R
XU11 VSS VDD  n6 n5 Output[2] XOR2xp5_ASAP7_75t_R
XU12 VSS VDD  n7 n8 INVx1_ASAP7_75t_R
XU13 VSS VDD  B[2] A[2] n10 NAND2xp5_ASAP7_75t_R
XU14 VSS VDD  n8 n10 n14 NAND2xp5_ASAP7_75t_R
XU15 VSS VDD  B[2] A[2] n13 OR2x2_ASAP7_75t_R
XU16 VSS VDD  n11 n10 n9 n12 NAND3xp33_ASAP7_75t_R
XU17 VSS VDD  n14 n13 n12 n16 NAND3xp33_ASAP7_75t_R
XU18 VSS VDD  B[3] A[3] n15 XNOR2xp5_ASAP7_75t_R
XU19 VSS VDD  n16 n15 Output[3] XOR2xp5_ASAP7_75t_R
XU20 VSS VDD  n16 n18 INVx1_ASAP7_75t_R
XU21 VSS VDD  B[3] A[3] n17 OR2x2_ASAP7_75t_R
XU22 VSS VDD  n18 n17 n20 NAND2xp5_ASAP7_75t_R
XU23 VSS VDD  B[3] A[3] n19 NAND2xp5_ASAP7_75t_R
XU24 VSS VDD  n20 n19 Output[4] NAND2xp5_ASAP7_75t_R
.ENDS



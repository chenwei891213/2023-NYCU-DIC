.SUBCKT Convolution VSS VDD  IFM_0[3] IFM_0[2] IFM_0[1] IFM_0[0] IFM_1[3] IFM_1[2] IFM_1[1] IFM_1[0] IFM_2[3] IFM_2[2] IFM_2[1] IFM_2[0] IFM_3[3] IFM_3[2] IFM_3[1] IFM_3[0] INW_0[3] INW_0[2] INW_0[1] INW_0[0] INW_1[3] INW_1[2] INW_1[1] INW_1[0] INW_2[3] INW_2[2] INW_2[1] INW_2[0] INW_3[3] INW_3[2] INW_3[1] INW_3[0] Output[9] Output[8] Output[7] Output[6] Output[5] Output[4] Output[3] Output[2] Output[1] Output[0] 
Xmult_19 VSS VDD  IFM_0[3] IFM_0[2] IFM_0[1] IFM_0[0] INW_0[3] INW_0[2] INW_0[1] INW_0[0] N7 N6 N5 N4 N3 N2 N1 N0 Convolution_DW_mult_uns_3
Xmult_19_2 VSS VDD  IFM_1[3] IFM_1[2] IFM_1[1] IFM_1[0] INW_1[3] INW_1[2] INW_1[1] INW_1[0] N15 N14 N13 N12 N11 N10 N9 N8 Convolution_DW_mult_uns_2
Xmult_19_3 VSS VDD  IFM_2[3] IFM_2[2] IFM_2[1] IFM_2[0] INW_2[3] INW_2[2] INW_2[1] INW_2[0] N32 N31 N30 N29 N28 N27 N26 N25 Convolution_DW_mult_uns_1
Xmult_19_4 VSS VDD  IFM_3[3] IFM_3[2] IFM_3[1] IFM_3[0] INW_3[3] INW_3[2] INW_3[1] INW_3[0] N50 N49 N48 N47 N46 N45 N44 N43 Convolution_DW_mult_uns_0
Xadd_1_root_add_0_root_add_19_3 VSS VDD  N42 N42 N15 N14 N13 N12 N11 N10 N9 N8 N42 N42 N50 N49 N48 N47 N46 N45 N44 N43 N42 SYNOPSYS_UNCONNECTED_1 new9 new8 new7 new6 new5 new4 new3 new2 new1 Convolution_DW01_add_2
Xadd_2_root_add_0_root_add_19_3 VSS VDD  N42 N42 N7 N6 N5 N4 N3 N2 N1 N0 N42 N42 N32 N31 N30 N29 N28 N27 N26 N25 N42 SYNOPSYS_UNCONNECTED_2 N41 N40 N39 N38 N37 N36 N35 N34 N33 Convolution_DW01_add_1
Xadd_0_root_add_0_root_add_19_3 VSS VDD  N42 N41 N40 N39 N38 N37 N36 N35 N34 N33 N42 new9 new8 new7 new6 new5 new4 new3 new2 new1 N42 Output[9] Output[8] Output[7] Output[6] Output[5] Output[4] Output[3] Output[2] Output[1] Output[0] Convolution_DW01_add_0
XU1 VSS VDD  N42 TIELOx1_ASAP7_75t_R
.ENDS


.SUBCKT  Convolution_DW01_add_0 VSS VDD A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] B[9] B[8] B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] CI SUM[9] SUM[8] SUM[7] SUM[6] SUM[5] SUM[4] SUM[3] SUM[2] SUM[1] SUM[0] 
XU1_8 VSS VDD  A[8] B[8] newa3 newa10 newa11 FAx1_ASAP7_75t_R
XU1_7 VSS VDD  A[7] B[7] newa4 newa12 newa13 FAx1_ASAP7_75t_R
XU1_6 VSS VDD  A[6] B[6] newa5 newa14 newa15 FAx1_ASAP7_75t_R
XU1_5 VSS VDD  A[5] B[5] newa6 newa16 newa17 FAx1_ASAP7_75t_R
XU1_4 VSS VDD  A[4] B[4] newa7 newa18 newa19 FAx1_ASAP7_75t_R
XU1_3 VSS VDD  A[3] B[3] newa8 newa20 newa21 FAx1_ASAP7_75t_R
XU1_2 VSS VDD  A[2] B[2] newa9 newa22 newa23 FAx1_ASAP7_75t_R
XU1_1 VSS VDD  A[1] B[1] newa1 newa24 newa25 FAx1_ASAP7_75t_R
XU1 VSS VDD  A[0] B[0] newa1 AND2x2_ASAP7_75t_R
XU2 VSS VDD  B[0] A[0] SUM[0] XOR2xp5_ASAP7_75t_R
XU3 VSS VDD  newa12 newa3 INVx1_ASAP7_75t_R
XU4 VSS VDD  newa14 newa4 INVx1_ASAP7_75t_R
XU5 VSS VDD  newa16 newa5 INVx1_ASAP7_75t_R
XU6 VSS VDD  newa18 newa6 INVx1_ASAP7_75t_R
XU7 VSS VDD  newa20 newa7 INVx1_ASAP7_75t_R
XU8 VSS VDD  newa22 newa8 INVx1_ASAP7_75t_R
XU9 VSS VDD  newa24 newa9 INVx1_ASAP7_75t_R
XU10 VSS VDD  newa10 SUM[9] INVx1_ASAP7_75t_R
XU11 VSS VDD  newa11 SUM[8] INVx1_ASAP7_75t_R
XU12 VSS VDD  newa13 SUM[7] INVx1_ASAP7_75t_R
XU13 VSS VDD  newa15 SUM[6] INVx1_ASAP7_75t_R
XU14 VSS VDD  newa17 SUM[5] INVx1_ASAP7_75t_R
XU15 VSS VDD  newa19 SUM[4] INVx1_ASAP7_75t_R
XU16 VSS VDD  newa21 SUM[3] INVx1_ASAP7_75t_R
XU17 VSS VDD  newa23 SUM[2] INVx1_ASAP7_75t_R
XU18 VSS VDD  newa25 SUM[1] INVx1_ASAP7_75t_R
.ENDS


.SUBCKT Convolution_DW01_add_1  VSS VDD A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] B[9] B[8] B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] CI SUM[9] SUM[8] SUM[7] SUM[6] SUM[5] SUM[4] SUM[3] SUM[2] SUM[1] SUM[0] 
XU1_7 VSS VDD  A[7] B[7] newb3 newb9 newb10 FAx1_ASAP7_75t_R
XU1_6 VSS VDD  A[6] B[6] newb4 newb11 newb12 FAx1_ASAP7_75t_R
XU1_5 VSS VDD  A[5] B[5] newb5 newb13 newb14 FAx1_ASAP7_75t_R
XU1_4 VSS VDD  A[4] B[4] newb6 newb15 newb16 FAx1_ASAP7_75t_R
XU1_3 VSS VDD  A[3] B[3] newb7 newb17 newb18 FAx1_ASAP7_75t_R
XU1_2 VSS VDD  A[2] B[2] newb8 newb19 newb20 FAx1_ASAP7_75t_R
XU1_1 VSS VDD  A[1] B[1] newb2 newb21 newb22 FAx1_ASAP7_75t_R
XU1 VSS VDD  B[0] A[0] SUM[0] XOR2xp5_ASAP7_75t_R
XU2 VSS VDD  A[0] B[0] newb2 AND2x2_ASAP7_75t_R
XU3 VSS VDD  newb11 newb3 INVx1_ASAP7_75t_R
XU4 VSS VDD  newb13 newb4 INVx1_ASAP7_75t_R
XU5 VSS VDD  newb15 newb5 INVx1_ASAP7_75t_R
XU6 VSS VDD  newb17 newb6 INVx1_ASAP7_75t_R
XU7 VSS VDD  newb19 newb7 INVx1_ASAP7_75t_R
XU8 VSS VDD  newb21 newb8 INVx1_ASAP7_75t_R
XU9 VSS VDD  newb9 SUM[8] INVx1_ASAP7_75t_R
XU10 VSS VDD  newb10 SUM[7] INVx1_ASAP7_75t_R
XU11 VSS VDD  newb12 SUM[6] INVx1_ASAP7_75t_R
XU12 VSS VDD  newb14 SUM[5] INVx1_ASAP7_75t_R
XU13 VSS VDD  newb16 SUM[4] INVx1_ASAP7_75t_R
XU14 VSS VDD  newb18 SUM[3] INVx1_ASAP7_75t_R
XU15 VSS VDD  newb20 SUM[2] INVx1_ASAP7_75t_R
XU16 VSS VDD  newb22 SUM[1] INVx1_ASAP7_75t_R
.ENDS


.SUBCKT  Convolution_DW01_add_2 VSS VDD A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] B[9] B[8] B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] CI SUM[9] SUM[8] SUM[7] SUM[6] SUM[5] SUM[4] SUM[3] SUM[2] SUM[1] SUM[0] 
XU1_7 VSS VDD  A[7] B[7] newc3 newc9 newc10 FAx1_ASAP7_75t_R
XU1_6 VSS VDD  A[6] B[6] newc4 newc11 newc12 FAx1_ASAP7_75t_R
XU1_5 VSS VDD  A[5] B[5] newc5 newc13 newc14 FAx1_ASAP7_75t_R
XU1_4 VSS VDD  A[4] B[4] newc6 newc15 newc16 FAx1_ASAP7_75t_R
XU1_3 VSS VDD  A[3] B[3] newc7 newc17 newc18 FAx1_ASAP7_75t_R
XU1_2 VSS VDD  A[2] B[2] newc8 newc19 newc20 FAx1_ASAP7_75t_R
XU1_1 VSS VDD  A[1] B[1] newc1 newc21 newc22 FAx1_ASAP7_75t_R
XU1 VSS VDD  A[0] B[0] newc1 AND2x2_ASAP7_75t_R
XU2 VSS VDD  B[0] A[0] SUM[0] XOR2xp5_ASAP7_75t_R
XU3 VSS VDD  newc11 newc3 INVx1_ASAP7_75t_R
XU4 VSS VDD  newc13 newc4 INVx1_ASAP7_75t_R
XU5 VSS VDD  newc15 newc5 INVx1_ASAP7_75t_R
XU6 VSS VDD  newc17 newc6 INVx1_ASAP7_75t_R
XU7 VSS VDD  newc19 newc7 INVx1_ASAP7_75t_R
XU8 VSS VDD  newc21 newc8 INVx1_ASAP7_75t_R
XU9 VSS VDD  newc9 SUM[8] INVx1_ASAP7_75t_R
XU10 VSS VDD  newc10 SUM[7] INVx1_ASAP7_75t_R
XU11 VSS VDD  newc12 SUM[6] INVx1_ASAP7_75t_R
XU12 VSS VDD  newc14 SUM[5] INVx1_ASAP7_75t_R
XU13 VSS VDD  newc16 SUM[4] INVx1_ASAP7_75t_R
XU14 VSS VDD  newc18 SUM[3] INVx1_ASAP7_75t_R
XU15 VSS VDD  newc20 SUM[2] INVx1_ASAP7_75t_R
XU16 VSS VDD  newc22 SUM[1] INVx1_ASAP7_75t_R
.ENDS


.SUBCKT  Convolution_DW_mult_uns_0 VSS VDD a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 VSS VDD  newd41 newd44 newd31 newd25 newd26 FAx1_ASAP7_75t_R
XU35 VSS VDD  newd36 newd45 newd32 newd29 newd30 FAx1_ASAP7_75t_R
XU39 VSS VDD  newd49 newd52 newd38 newd34 newd35 FAx1_ASAP7_75t_R
XU70 VSS VDD  a[2] newd83 INVx1_ASAP7_75t_R
XU71 VSS VDD  newd35 newd84 INVx1_ASAP7_75t_R
XU72 VSS VDD  a[0] newd85 INVx1_ASAP7_75t_R
XU73 VSS VDD  b[3] newd86 INVx1_ASAP7_75t_R
XU74 VSS VDD  b[0] newd87 INVx1_ASAP7_75t_R
XU75 VSS VDD  newd88 newd89 product[7] NAND2xp33_ASAP7_75t_R
XU76 VSS VDD  newd90 newd91 newd89 NAND2xp33_ASAP7_75t_R
XU77 VSS VDD  newd92 newd25 newd88 OR2x2_ASAP7_75t_R
XU78 VSS VDD  newd91 newd90 product[6] XOR2xp5_ASAP7_75t_R
XU79 VSS VDD  newd92 newd25 newd90 XOR2xp5_ASAP7_75t_R
XU80 VSS VDD  b[3] a[3] newd92 NAND2xp33_ASAP7_75t_R
XU81 VSS VDD  newd93 newd94 newd91 NAND2xp33_ASAP7_75t_R
XU82 VSS VDD  newd95 newd96 newd94 NAND2xp33_ASAP7_75t_R
XU83 VSS VDD  newd26 newd29 newd93 OR2x2_ASAP7_75t_R
XU84 VSS VDD  newd96 newd95 product[5] XOR2xp5_ASAP7_75t_R
XU85 VSS VDD  newd26 newd29 newd95 XOR2xp5_ASAP7_75t_R
XU86 VSS VDD  newd97 newd98 newd96 NAND2xp33_ASAP7_75t_R
XU87 VSS VDD  newd99 newd100 newd98 NAND2xp33_ASAP7_75t_R
XU88 VSS VDD  newd30 newd34 newd97 OR2x2_ASAP7_75t_R
XU89 VSS VDD  newd100 newd99 product[4] XOR2xp5_ASAP7_75t_R
XU90 VSS VDD  newd30 newd34 newd99 XOR2xp5_ASAP7_75t_R
XU91 VSS VDD  newd101 newd102 newd100 NAND2xp33_ASAP7_75t_R
XU92 VSS VDD  newd103 newd104 newd102 NAND2xp33_ASAP7_75t_R
XU93 VSS VDD  newd105 newd84 newd101 NAND2xp33_ASAP7_75t_R
XU94 VSS VDD  newd104 newd103 product[3] XOR2xp5_ASAP7_75t_R
XU95 VSS VDD  newd35 newd105 newd103 XNOR2xp5_ASAP7_75t_R
XU96 VSS VDD  newd106 newd107 newd105 XOR2xp5_ASAP7_75t_R
XU97 VSS VDD  newd108 newd109 newd104 NAND2xp33_ASAP7_75t_R
XU98 VSS VDD  newd110 newd111 newd109 NAND2xp33_ASAP7_75t_R
XU99 VSS VDD  newd112 newd113 newd108 NAND2xp33_ASAP7_75t_R
XU100 VSS VDD  newd110 newd111 product[2] XOR2xp5_ASAP7_75t_R
XU101 VSS VDD  newd112 newd113 newd111 XOR2xp5_ASAP7_75t_R
XU102 VSS VDD  newd114 newd115 newd113 XOR2xp5_ASAP7_75t_R
XU103 VSS VDD  newd83 newd87 newd112 NOR2xp33_ASAP7_75t_R
XU104 VSS VDD  newd116 newd117 newd110 NOR2xp33_ASAP7_75t_R
XU105 VSS VDD  newd116 newd117 product[1] XOR2xp5_ASAP7_75t_R
XU106 VSS VDD  b[1] a[0] newd117 NAND2xp33_ASAP7_75t_R
XU107 VSS VDD  b[0] a[1] newd116 NAND2xp33_ASAP7_75t_R
XU108 VSS VDD  newd87 newd85 product[0] NOR2xp33_ASAP7_75t_R
XU109 VSS VDD  newd85 newd86 newd52 NOR2xp33_ASAP7_75t_R
XU110 VSS VDD  a[1] b[2] newd49 AND2x2_ASAP7_75t_R
XU111 VSS VDD  a[2] b[2] newd45 AND2x2_ASAP7_75t_R
XU112 VSS VDD  newd83 newd86 newd44 NOR2xp33_ASAP7_75t_R
XU113 VSS VDD  b[2] a[3] newd41 AND2x2_ASAP7_75t_R
XU114 VSS VDD  newd115 newd114 newd38 NOR2xp33_ASAP7_75t_R
XU115 VSS VDD  b[1] a[1] newd114 NAND2xp33_ASAP7_75t_R
XU116 VSS VDD  b[2] a[0] newd115 NAND2xp33_ASAP7_75t_R
XU117 VSS VDD  newd107 newd106 newd36 NOR2xp33_ASAP7_75t_R
XU118 VSS VDD  a[3] b[0] newd106 NAND2xp33_ASAP7_75t_R
XU119 VSS VDD  a[2] b[1] newd107 NAND2xp33_ASAP7_75t_R
XU120 VSS VDD  newd118 newd119 newd32 XOR2xp5_ASAP7_75t_R
XU121 VSS VDD  newd118 newd119 newd31 NOR2xp33_ASAP7_75t_R
XU122 VSS VDD  a[3] b[1] newd119 NAND2xp33_ASAP7_75t_R
XU123 VSS VDD  b[3] a[1] newd118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT  Convolution_DW_mult_uns_1 VSS VDD a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 VSS VDD  newe41 newe44 newe31 newe25 newe26 FAx1_ASAP7_75t_R
XU35 VSS VDD  newe36 newe45 newe32 newe29 newe30 FAx1_ASAP7_75t_R
XU39 VSS VDD  newe49 newe52 newe38 newe34 newe35 FAx1_ASAP7_75t_R
XU70 VSS VDD  a[2] newe83 INVx1_ASAP7_75t_R
XU71 VSS VDD  newe35 newe84 INVx1_ASAP7_75t_R
XU72 VSS VDD  a[0] newe85 INVx1_ASAP7_75t_R
XU73 VSS VDD  b[3] newe86 INVx1_ASAP7_75t_R
XU74 VSS VDD  b[0] newe87 INVx1_ASAP7_75t_R
XU75 VSS VDD  newe88 newe89 product[7] NAND2xp33_ASAP7_75t_R
XU76 VSS VDD  newe90 newe91 newe89 NAND2xp33_ASAP7_75t_R
XU77 VSS VDD  newe92 newe25 newe88 OR2x2_ASAP7_75t_R
XU78 VSS VDD  newe91 newe90 product[6] XOR2xp5_ASAP7_75t_R
XU79 VSS VDD  newe92 newe25 newe90 XOR2xp5_ASAP7_75t_R
XU80 VSS VDD  b[3] a[3] newe92 NAND2xp33_ASAP7_75t_R
XU81 VSS VDD  newe93 newe94 newe91 NAND2xp33_ASAP7_75t_R
XU82 VSS VDD  newe95 newe96 newe94 NAND2xp33_ASAP7_75t_R
XU83 VSS VDD  newe26 newe29 newe93 OR2x2_ASAP7_75t_R
XU84 VSS VDD  newe96 newe95 product[5] XOR2xp5_ASAP7_75t_R
XU85 VSS VDD  newe26 newe29 newe95 XOR2xp5_ASAP7_75t_R
XU86 VSS VDD  newe97 newe98 newe96 NAND2xp33_ASAP7_75t_R
XU87 VSS VDD  newe99 newe100 newe98 NAND2xp33_ASAP7_75t_R
XU88 VSS VDD  newe30 newe34 newe97 OR2x2_ASAP7_75t_R
XU89 VSS VDD  newe100 newe99 product[4] XOR2xp5_ASAP7_75t_R
XU90 VSS VDD  newe30 newe34 newe99 XOR2xp5_ASAP7_75t_R
XU91 VSS VDD  newe101 newe102 newe100 NAND2xp33_ASAP7_75t_R
XU92 VSS VDD  newe103 newe104 newe102 NAND2xp33_ASAP7_75t_R
XU93 VSS VDD  newe105 newe84 newe101 NAND2xp33_ASAP7_75t_R
XU94 VSS VDD  newe104 newe103 product[3] XOR2xp5_ASAP7_75t_R
XU95 VSS VDD  newe35 newe105 newe103 XNOR2xp5_ASAP7_75t_R
XU96 VSS VDD  newe106 newe107 newe105 XOR2xp5_ASAP7_75t_R
XU97 VSS VDD  newe108 newe109 newe104 NAND2xp33_ASAP7_75t_R
XU98 VSS VDD  newe110 newe111 newe109 NAND2xp33_ASAP7_75t_R
XU99 VSS VDD  newe112 newe113 newe108 NAND2xp33_ASAP7_75t_R
XU100 VSS VDD  newe110 newe111 product[2] XOR2xp5_ASAP7_75t_R
XU101 VSS VDD  newe112 newe113 newe111 XOR2xp5_ASAP7_75t_R
XU102 VSS VDD  newe114 newe115 newe113 XOR2xp5_ASAP7_75t_R
XU103 VSS VDD  newe83 newe87 newe112 NOR2xp33_ASAP7_75t_R
XU104 VSS VDD  newe116 newe117 newe110 NOR2xp33_ASAP7_75t_R
XU105 VSS VDD  newe116 newe117 product[1] XOR2xp5_ASAP7_75t_R
XU106 VSS VDD  b[1] a[0] newe117 NAND2xp33_ASAP7_75t_R
XU107 VSS VDD  b[0] a[1] newe116 NAND2xp33_ASAP7_75t_R
XU108 VSS VDD  newe87 newe85 product[0] NOR2xp33_ASAP7_75t_R
XU109 VSS VDD  newe85 newe86 newe52 NOR2xp33_ASAP7_75t_R
XU110 VSS VDD  a[1] b[2] newe49 AND2x2_ASAP7_75t_R
XU111 VSS VDD  a[2] b[2] newe45 AND2x2_ASAP7_75t_R
XU112 VSS VDD  newe83 newe86 newe44 NOR2xp33_ASAP7_75t_R
XU113 VSS VDD  b[2] a[3] newe41 AND2x2_ASAP7_75t_R
XU114 VSS VDD  newe115 newe114 newe38 NOR2xp33_ASAP7_75t_R
XU115 VSS VDD  b[1] a[1] newe114 NAND2xp33_ASAP7_75t_R
XU116 VSS VDD  b[2] a[0] newe115 NAND2xp33_ASAP7_75t_R
XU117 VSS VDD  newe107 newe106 newe36 NOR2xp33_ASAP7_75t_R
XU118 VSS VDD  a[3] b[0] newe106 NAND2xp33_ASAP7_75t_R
XU119 VSS VDD  a[2] b[1] newe107 NAND2xp33_ASAP7_75t_R
XU120 VSS VDD  newe118 newe119 newe32 XOR2xp5_ASAP7_75t_R
XU121 VSS VDD  newe118 newe119 newe31 NOR2xp33_ASAP7_75t_R
XU122 VSS VDD  a[3] b[1] newe119 NAND2xp33_ASAP7_75t_R
XU123 VSS VDD  b[3] a[1] newe118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT Convolution_DW_mult_uns_2  VSS VDD a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 VSS VDD  newf41 newf44 newf31 newf25 newf26 FAx1_ASAP7_75t_R
XU35 VSS VDD  newf36 newf45 newf32 newf29 newf30 FAx1_ASAP7_75t_R
XU39 VSS VDD  newf49 newf52 newf38 newf34 newf35 FAx1_ASAP7_75t_R
XU70 VSS VDD  a[2] newf83 INVx1_ASAP7_75t_R
XU71 VSS VDD  newf35 newf84 INVx1_ASAP7_75t_R
XU72 VSS VDD  a[0] newf85 INVx1_ASAP7_75t_R
XU73 VSS VDD  b[3] newf86 INVx1_ASAP7_75t_R
XU74 VSS VDD  b[0] newf87 INVx1_ASAP7_75t_R
XU75 VSS VDD  newf88 newf89 product[7] NAND2xp33_ASAP7_75t_R
XU76 VSS VDD  newf90 newf91 newf89 NAND2xp33_ASAP7_75t_R
XU77 VSS VDD  newf92 newf25 newf88 OR2x2_ASAP7_75t_R
XU78 VSS VDD  newf91 newf90 product[6] XOR2xp5_ASAP7_75t_R
XU79 VSS VDD  newf92 newf25 newf90 XOR2xp5_ASAP7_75t_R
XU80 VSS VDD  b[3] a[3] newf92 NAND2xp33_ASAP7_75t_R
XU81 VSS VDD  newf93 newf94 newf91 NAND2xp33_ASAP7_75t_R
XU82 VSS VDD  newf95 newf96 newf94 NAND2xp33_ASAP7_75t_R
XU83 VSS VDD  newf26 newf29 newf93 OR2x2_ASAP7_75t_R
XU84 VSS VDD  newf96 newf95 product[5] XOR2xp5_ASAP7_75t_R
XU85 VSS VDD  newf26 newf29 newf95 XOR2xp5_ASAP7_75t_R
XU86 VSS VDD  newf97 newf98 newf96 NAND2xp33_ASAP7_75t_R
XU87 VSS VDD  newf99 newf100 newf98 NAND2xp33_ASAP7_75t_R
XU88 VSS VDD  newf30 newf34 newf97 OR2x2_ASAP7_75t_R
XU89 VSS VDD  newf100 newf99 product[4] XOR2xp5_ASAP7_75t_R
XU90 VSS VDD  newf30 newf34 newf99 XOR2xp5_ASAP7_75t_R
XU91 VSS VDD  newf101 newf102 newf100 NAND2xp33_ASAP7_75t_R
XU92 VSS VDD  newf103 newf104 newf102 NAND2xp33_ASAP7_75t_R
XU93 VSS VDD  newf105 newf84 newf101 NAND2xp33_ASAP7_75t_R
XU94 VSS VDD  newf104 newf103 product[3] XOR2xp5_ASAP7_75t_R
XU95 VSS VDD  newf35 newf105 newf103 XNOR2xp5_ASAP7_75t_R
XU96 VSS VDD  newf106 newf107 newf105 XOR2xp5_ASAP7_75t_R
XU97 VSS VDD  newf108 newf109 newf104 NAND2xp33_ASAP7_75t_R
XU98 VSS VDD  newf110 newf111 newf109 NAND2xp33_ASAP7_75t_R
XU99 VSS VDD  newf112 newf113 newf108 NAND2xp33_ASAP7_75t_R
XU100 VSS VDD  newf110 newf111 product[2] XOR2xp5_ASAP7_75t_R
XU101 VSS VDD  newf112 newf113 newf111 XOR2xp5_ASAP7_75t_R
XU102 VSS VDD  newf114 newf115 newf113 XOR2xp5_ASAP7_75t_R
XU103 VSS VDD  newf83 newf87 newf112 NOR2xp33_ASAP7_75t_R
XU104 VSS VDD  newf116 newf117 newf110 NOR2xp33_ASAP7_75t_R
XU105 VSS VDD  newf116 newf117 product[1] XOR2xp5_ASAP7_75t_R
XU106 VSS VDD  b[1] a[0] newf117 NAND2xp33_ASAP7_75t_R
XU107 VSS VDD  b[0] a[1] newf116 NAND2xp33_ASAP7_75t_R
XU108 VSS VDD  newf87 newf85 product[0] NOR2xp33_ASAP7_75t_R
XU109 VSS VDD  newf85 newf86 newf52 NOR2xp33_ASAP7_75t_R
XU110 VSS VDD  a[1] b[2] newf49 AND2x2_ASAP7_75t_R
XU111 VSS VDD  a[2] b[2] newf45 AND2x2_ASAP7_75t_R
XU112 VSS VDD  newf83 newf86 newf44 NOR2xp33_ASAP7_75t_R
XU113 VSS VDD  b[2] a[3] newf41 AND2x2_ASAP7_75t_R
XU114 VSS VDD  newf115 newf114 newf38 NOR2xp33_ASAP7_75t_R
XU115 VSS VDD  b[1] a[1] newf114 NAND2xp33_ASAP7_75t_R
XU116 VSS VDD  b[2] a[0] newf115 NAND2xp33_ASAP7_75t_R
XU117 VSS VDD  newf107 newf106 newf36 NOR2xp33_ASAP7_75t_R
XU118 VSS VDD  a[3] b[0] newf106 NAND2xp33_ASAP7_75t_R
XU119 VSS VDD  a[2] b[1] newf107 NAND2xp33_ASAP7_75t_R
XU120 VSS VDD  newf118 newf119 newf32 XOR2xp5_ASAP7_75t_R
XU121 VSS VDD  newf118 newf119 newf31 NOR2xp33_ASAP7_75t_R
XU122 VSS VDD  a[3] b[1] newf119 NAND2xp33_ASAP7_75t_R
XU123 VSS VDD  b[3] a[1] newf118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT Convolution_DW_mult_uns_3 VSS VDD  a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 VSS VDD  newg41 newg44 newg31 newg25 newg26 FAx1_ASAP7_75t_R
XU35 VSS VDD  newg36 newg45 newg32 newg29 newg30 FAx1_ASAP7_75t_R
XU39 VSS VDD  newg49 newg52 newg38 newg34 newg35 FAx1_ASAP7_75t_R
XU70 VSS VDD  a[2] newg83 INVx1_ASAP7_75t_R
XU71 VSS VDD  newg35 newg84 INVx1_ASAP7_75t_R
XU72 VSS VDD  a[0] newg85 INVx1_ASAP7_75t_R
XU73 VSS VDD  b[3] newg86 INVx1_ASAP7_75t_R
XU74 VSS VDD  b[0] newg87 INVx1_ASAP7_75t_R
XU75 VSS VDD  newg88 newg89 product[7] NAND2xp33_ASAP7_75t_R
XU76 VSS VDD  newg90 newg91 newg89 NAND2xp33_ASAP7_75t_R
XU77 VSS VDD  newg92 newg25 newg88 OR2x2_ASAP7_75t_R
XU78 VSS VDD  newg91 newg90 product[6] XOR2xp5_ASAP7_75t_R
XU79 VSS VDD  newg92 newg25 newg90 XOR2xp5_ASAP7_75t_R
XU80 VSS VDD  b[3] a[3] newg92 NAND2xp33_ASAP7_75t_R
XU81 VSS VDD  newg93 newg94 newg91 NAND2xp33_ASAP7_75t_R
XU82 VSS VDD  newg95 newg96 newg94 NAND2xp33_ASAP7_75t_R
XU83 VSS VDD  newg26 newg29 newg93 OR2x2_ASAP7_75t_R
XU84 VSS VDD  newg96 newg95 product[5] XOR2xp5_ASAP7_75t_R
XU85 VSS VDD  newg26 newg29 newg95 XOR2xp5_ASAP7_75t_R
XU86 VSS VDD  newg97 newg98 newg96 NAND2xp33_ASAP7_75t_R
XU87 VSS VDD  newg99 newg100 newg98 NAND2xp33_ASAP7_75t_R
XU88 VSS VDD  newg30 newg34 newg97 OR2x2_ASAP7_75t_R
XU89 VSS VDD  newg100 newg99 product[4] XOR2xp5_ASAP7_75t_R
XU90 VSS VDD  newg30 newg34 newg99 XOR2xp5_ASAP7_75t_R
XU91 VSS VDD  newg101 newg102 newg100 NAND2xp33_ASAP7_75t_R
XU92 VSS VDD  newg103 newg104 newg102 NAND2xp33_ASAP7_75t_R
XU93 VSS VDD  newg105 newg84 newg101 NAND2xp33_ASAP7_75t_R
XU94 VSS VDD  newg104 newg103 product[3] XOR2xp5_ASAP7_75t_R
XU95 VSS VDD  newg35 newg105 newg103 XNOR2xp5_ASAP7_75t_R
XU96 VSS VDD  newg106 newg107 newg105 XOR2xp5_ASAP7_75t_R
XU97 VSS VDD  newg108 newg109 newg104 NAND2xp33_ASAP7_75t_R
XU98 VSS VDD  newg110 newg111 newg109 NAND2xp33_ASAP7_75t_R
XU99 VSS VDD  newg112 newg113 newg108 NAND2xp33_ASAP7_75t_R
XU100 VSS VDD  newg110 newg111 product[2] XOR2xp5_ASAP7_75t_R
XU101 VSS VDD  newg112 newg113 newg111 XOR2xp5_ASAP7_75t_R
XU102 VSS VDD  newg114 newg115 newg113 XOR2xp5_ASAP7_75t_R
XU103 VSS VDD  newg83 newg87 newg112 NOR2xp33_ASAP7_75t_R
XU104 VSS VDD  newg116 newg117 newg110 NOR2xp33_ASAP7_75t_R
XU105 VSS VDD  newg116 newg117 product[1] XOR2xp5_ASAP7_75t_R
XU106 VSS VDD  b[1] a[0] newg117 NAND2xp33_ASAP7_75t_R
XU107 VSS VDD  b[0] a[1] newg116 NAND2xp33_ASAP7_75t_R
XU108 VSS VDD  newg87 newg85 product[0] NOR2xp33_ASAP7_75t_R
XU109 VSS VDD  newg85 newg86 newg52 NOR2xp33_ASAP7_75t_R
XU110 VSS VDD  a[1] b[2] newg49 AND2x2_ASAP7_75t_R
XU111 VSS VDD  a[2] b[2] newg45 AND2x2_ASAP7_75t_R
XU112 VSS VDD  newg83 newg86 newg44 NOR2xp33_ASAP7_75t_R
XU113 VSS VDD  b[2] a[3] newg41 AND2x2_ASAP7_75t_R
XU114 VSS VDD  newg115 newg114 newg38 NOR2xp33_ASAP7_75t_R
XU115 VSS VDD  b[1] a[1] newg114 NAND2xp33_ASAP7_75t_R
XU116 VSS VDD  b[2] a[0] newg115 NAND2xp33_ASAP7_75t_R
XU117 VSS VDD  newg107 newg106 newg36 NOR2xp33_ASAP7_75t_R
XU118 VSS VDD  a[3] b[0] newg106 NAND2xp33_ASAP7_75t_R
XU119 VSS VDD  a[2] b[1] newg107 NAND2xp33_ASAP7_75t_R
XU120 VSS VDD  newg118 newg119 newg32 XOR2xp5_ASAP7_75t_R
XU121 VSS VDD  newg118 newg119 newg31 NOR2xp33_ASAP7_75t_R
XU122 VSS VDD  a[3] b[1] newg119 NAND2xp33_ASAP7_75t_R
XU123 VSS VDD  b[3] a[1] newg118 NAND2xp33_ASAP7_75t_R
.ENDS



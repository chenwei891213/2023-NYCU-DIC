* Design:	DFFHQNx1_ASAP7_75t_R
* Created:	"Fri Aug 17 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "DFFHQNx1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "DFFHQNx1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_DFFHQNx1_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.00427064f
.ends

.subckt PM_DFFHQNx1_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.00416001f
.ends

.subckt PM_DFFHQNx1_ASAP7_75t_R%noxref_29 VSS 1
c1 1 VSS 0.00452737f
.ends

.subckt PM_DFFHQNx1_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.00426212f
.ends

.subckt PM_DFFHQNx1_ASAP7_75t_R%noxref_28 VSS 1
c1 1 VSS 0.00477846f
.ends

.subckt PM_DFFHQNx1_ASAP7_75t_R%noxref_26 VSS 1
c1 1 VSS 0.0415028f
.ends

.subckt PM_DFFHQNx1_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.00426485f
.ends

.subckt PM_DFFHQNx1_ASAP7_75t_R%noxref_27 VSS 1
c1 1 VSS 0.0415009f
.ends

.subckt PM_DFFHQNx1_ASAP7_75t_R%QN VSS 19 13 25 2 7 9 1 8
c1 1 VSS 0.00826277f
c2 2 VSS 0.00838008f
c3 7 VSS 0.00367384f
c4 8 VSS 0.00366397f
c5 9 VSS 0.00332205f
c6 10 VSS 0.00624757f
c7 11 VSS 0.00582331f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0115 $Y=0.2025 $X2=1.0240 $Y2=0.2025
r2 25 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0090 $Y=0.2025 $X2=1.0115 $Y2=0.2025
r3 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0260 $Y=0.2025
+ $X2=1.0260 $Y2=0.2340
r4 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.2340 $X2=1.0395 $Y2=0.2340
r5 11 20 1.09329 $w=1.76154e-08 $l=9.8e-09 $layer=M1 $thickness=3.6e-08
+ $X=1.0530 $Y=0.2340 $X2=1.0530 $Y2=0.2242
r6 11 23 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0530 $Y=0.2340 $X2=1.0395 $Y2=0.2340
r7 19 20 0.291487 $w=1.3e-08 $l=1.2e-09 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.2230 $X2=1.0530 $Y2=0.2242
r8 19 18 6.58761 $w=1.3e-08 $l=2.83e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.2230 $X2=1.0530 $Y2=0.1947
r9 17 18 15.4488 $w=1.3e-08 $l=6.62e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1285 $X2=1.0530 $Y2=0.1947
r10 9 16 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0530 $Y=0.0675 $X2=1.0530 $Y2=0.0360
r11 9 17 14.2246 $w=1.3e-08 $l=6.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.0675 $X2=1.0530 $Y2=0.1285
r12 15 16 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0395 $Y=0.0360 $X2=1.0530 $Y2=0.0360
r13 14 15 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.0360 $X2=1.0395 $Y2=0.0360
r14 10 14 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.0145
+ $Y=0.0360 $X2=1.0260 $Y2=0.0360
r15 1 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0260 $Y=0.0675
+ $X2=1.0260 $Y2=0.0360
r16 7 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.0115 $Y=0.0675 $X2=1.0240 $Y2=0.0675
r17 13 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.0090 $Y=0.0675 $X2=1.0115 $Y2=0.0675
.ends

.subckt PM_DFFHQNx1_ASAP7_75t_R%PD3 VSS 2 4 1
c1 1 VSS 0.000972222f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0405 $X2=0.4905 $Y2=0.0405
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0405 $X2=0.4735 $Y2=0.0405
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4735 $Y=0.0405 $X2=0.4905 $Y2=0.0405
.ends

.subckt PM_DFFHQNx1_ASAP7_75t_R%PD4 VSS 2 4 1
c1 1 VSS 0.000945784f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.2295 $X2=0.7605 $Y2=0.2295
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.2295 $X2=0.7435 $Y2=0.2295
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7435 $Y=0.2295 $X2=0.7605 $Y2=0.2295
.ends

.subckt PM_DFFHQNx1_ASAP7_75t_R%PU1 VSS 2 4 1
c1 1 VSS 0.0009845f
r1 4 3 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3365 $Y2=0.2025
r2 2 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3195 $Y2=0.2025
r3 1 3 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3195 $Y=0.2025 $X2=0.3365 $Y2=0.2025
.ends

.subckt PM_DFFHQNx1_ASAP7_75t_R%PD2 VSS 7 12 4 5 1
c1 1 VSS 0.00730038f
c2 4 VSS 0.00188731f
c3 5 VSS 0.00233441f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4880 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r3 9 5 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.4605
+ $Y=0.2295 $X2=0.4860 $Y2=0.2295
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.4455
+ $Y=0.2295 $X2=0.4605 $Y2=0.2295
r5 1 8 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4320
+ $Y=0.2295 $X2=0.4455 $Y2=0.2295
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2295 $X2=0.4300 $Y2=0.2295
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2295 $X2=0.4175 $Y2=0.2295
.ends

.subckt PM_DFFHQNx1_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.00485299f
.ends

.subckt PM_DFFHQNx1_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.041561f
.ends

.subckt PM_DFFHQNx1_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.00487019f
.ends

.subckt PM_DFFHQNx1_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.0415701f
.ends

.subckt PM_DFFHQNx1_ASAP7_75t_R%SS VSS 9 31 41 12 10 11 15 4 3 14 1 16 13 17
c1 1 VSS 0.00102999f
c2 3 VSS 0.00624336f
c3 4 VSS 0.00663106f
c4 9 VSS 0.0384397f
c5 10 VSS 0.00326083f
c6 11 VSS 0.00324511f
c7 12 VSS 0.00185534f
c8 13 VSS 0.0135942f
c9 14 VSS 0.00902919f
c10 15 VSS 0.00619638f
c11 16 VSS 0.00323914f
c12 17 VSS 0.00312957f
c13 18 VSS 0.00316281f
r1 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.2295 $X2=0.8620 $Y2=0.2295
r2 41 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.2295 $X2=0.8495 $Y2=0.2295
r3 4 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.2295
+ $X2=0.8640 $Y2=0.2340
r4 38 39 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.2340 $X2=0.8865 $Y2=0.2340
r5 14 18 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9180 $Y=0.2340 $X2=0.9450 $Y2=0.2340
r6 14 39 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.2340 $X2=0.8865 $Y2=0.2340
r7 18 36 0.56619 $w=2.22842e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.2340 $X2=0.9450 $Y2=0.2245
r8 35 36 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1975 $X2=0.9450 $Y2=0.2245
r9 34 35 6.64591 $w=1.3e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1690 $X2=0.9450 $Y2=0.1975
r10 33 34 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1420 $X2=0.9450 $Y2=0.1690
r11 32 33 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1035 $X2=0.9450 $Y2=0.1420
r12 15 17 5.69636 $w=1.58e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.0675 $X2=0.9450 $Y2=0.0360
r13 15 32 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.0675 $X2=0.9450 $Y2=0.1035
r14 10 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.0405 $X2=0.8620 $Y2=0.0405
r15 31 10 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.0405 $X2=0.8495 $Y2=0.0405
r16 17 29 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.0360 $X2=0.9180 $Y2=0.0360
r17 3 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.0405
+ $X2=0.8640 $Y2=0.0360
r18 28 29 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.0360 $X2=0.9180 $Y2=0.0360
r19 27 28 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.0360 $X2=0.8910 $Y2=0.0360
r20 26 27 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.0360 $X2=0.8640 $Y2=0.0360
r21 13 16 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.0360 $X2=0.7830 $Y2=0.0360
r22 13 26 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0360 $X2=0.8370 $Y2=0.0360
r23 12 23 8.04505 $w=1.3e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.0705 $X2=0.7830 $Y2=0.1050
r24 12 16 6.39593 $w=1.55565e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7830 $Y=0.0705 $X2=0.7830 $Y2=0.0360
r25 1 20 2.36633 $w=2.3e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.7830
+ $Y=0.1055 $X2=0.7830 $Y2=0.1055
r26 1 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7830 $Y=0.1055
+ $X2=0.7830 $Y2=0.1050
r27 9 20 0.314665 $w=2.27e-07 $l=2.95e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.7830 $Y=0.1350 $X2=0.7830 $Y2=0.1055
.ends

.subckt PM_DFFHQNx1_ASAP7_75t_R%PD5 VSS 7 12 4 1 5
c1 1 VSS 0.00741411f
c2 4 VSS 0.00187966f
c3 5 VSS 0.00237599f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.0405 $X2=0.7705 $Y2=0.0405
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7580 $Y=0.0405 $X2=0.7705 $Y2=0.0405
r3 9 5 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.7425
+ $Y=0.0405 $X2=0.7560 $Y2=0.0405
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.7275
+ $Y=0.0405 $X2=0.7425 $Y2=0.0405
r5 1 8 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.7020
+ $Y=0.0405 $X2=0.7275 $Y2=0.0405
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.0405 $X2=0.7000 $Y2=0.0405
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.0405 $X2=0.6875 $Y2=0.0405
.ends

.subckt PM_DFFHQNx1_ASAP7_75t_R%CLK VSS 10 3 8 5 1 6 7 4
c1 1 VSS 0.00247155f
c2 3 VSS 0.0596776f
c3 4 VSS 0.000945964f
c4 5 VSS 0.00399877f
c5 6 VSS 0.0038827f
c6 7 VSS 0.00219792f
c7 8 VSS 0.00206941f
r1 6 18 3.22357 $w=2.26279e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.2125 $X2=0.1080 $Y2=0.1820
r2 5 16 3.22357 $w=2.26279e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0575 $X2=0.1080 $Y2=0.0880
r3 17 18 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.1820 $X2=0.1080 $Y2=0.1820
r4 8 14 0.54189 $w=3.37e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1820 $X2=0.0810 $Y2=0.1630
r5 8 17 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1820 $X2=0.0945 $Y2=0.1820
r6 15 16 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.0880 $X2=0.1080 $Y2=0.0880
r7 7 15 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0880 $X2=0.0945 $Y2=0.0880
r8 13 14 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1530 $X2=0.0810 $Y2=0.1630
r9 12 13 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1530
r10 11 12 2.85657 $w=1.3e-08 $l=1.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1227 $X2=0.0810 $Y2=0.1350
r11 10 11 0.874462 $w=1.3e-08 $l=3.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1227
r12 10 4 1.57403 $w=1.3e-08 $l=6.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1122
r13 4 7 1.76614 $w=2.65738e-08 $l=2.42e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1122 $X2=0.0810 $Y2=0.0880
r14 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r15 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_DFFHQNx1_ASAP7_75t_R%MS VSS 10 41 44 48 50 13 17 18 14 3 15 12 1 11
+ 4 16
c1 1 VSS 0.00215722f
c2 3 VSS 0.00567637f
c3 4 VSS 0.0093574f
c4 10 VSS 0.0375163f
c5 11 VSS 0.00306316f
c6 12 VSS 0.00287648f
c7 13 VSS 0.00244325f
c8 14 VSS 0.00192209f
c9 15 VSS 0.00401872f
c10 16 VSS 0.00194786f
c11 17 VSS 0.0012613f
c12 18 VSS 0.000426788f
c13 19 VSS 0.00278384f
r1 50 49 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.2295 $X2=0.6625 $Y2=0.2295
r2 13 49 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6500 $Y=0.2295 $X2=0.6625 $Y2=0.2295
r3 12 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2295 $X2=0.5920 $Y2=0.2295
r4 48 12 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.2295 $X2=0.5795 $Y2=0.2295
r5 45 13 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6210 $Y=0.2295 $X2=0.6480 $Y2=0.2295
r6 4 45 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08 $X=0.5940
+ $Y=0.2295 $X2=0.6210 $Y2=0.2295
r7 4 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2295
+ $X2=0.5940 $Y2=0.2340
r8 15 19 5.06479 $w=1.46038e-08 $l=2.70046e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5940 $Y=0.2340 $X2=0.6210 $Y2=0.2335
r9 44 43 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.0405 $X2=0.6085 $Y2=0.0405
r10 42 43 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6040 $Y=0.0405 $X2=0.6085 $Y2=0.0405
r11 3 42 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5920 $Y=0.0405 $X2=0.6040 $Y2=0.0405
r12 11 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.0405 $X2=0.5920 $Y2=0.0405
r13 41 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0405 $X2=0.5795 $Y2=0.0405
r14 19 36 0.983973 $w=1.77222e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.2335 $X2=0.6210 $Y2=0.2245
r15 3 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0405
+ $X2=0.5940 $Y2=0.0540
r16 35 36 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.2135 $X2=0.6210 $Y2=0.2245
r17 34 35 6.64591 $w=1.3e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1850 $X2=0.6210 $Y2=0.2135
r18 33 34 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1660 $X2=0.6210 $Y2=0.1850
r19 32 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1525 $X2=0.6210 $Y2=0.1660
r20 31 32 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1310 $X2=0.6210 $Y2=0.1525
r21 30 31 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1115 $X2=0.6210 $Y2=0.1310
r22 17 28 1.15159 $w=1.75e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1000 $X2=0.6210 $Y2=0.0900
r23 17 30 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1000 $X2=0.6210 $Y2=0.1115
r24 16 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0540 $X2=0.5940 $Y2=0.0720
r25 27 28 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6075 $Y=0.0900 $X2=0.6210 $Y2=0.0900
r26 18 26 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5940 $Y=0.0900 $X2=0.5805 $Y2=0.0900
r27 18 27 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5940 $Y=0.0900 $X2=0.6075 $Y2=0.0900
r28 18 29 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0900 $X2=0.5940 $Y2=0.0720
r29 25 26 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5490
+ $Y=0.0900 $X2=0.5805 $Y2=0.0900
r30 24 25 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0900 $X2=0.5490 $Y2=0.0900
r31 14 24 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5000
+ $Y=0.0900 $X2=0.5130 $Y2=0.0900
r32 1 21 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.5130
+ $Y=0.0900 $X2=0.5130 $Y2=0.0900
r33 1 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.0900
+ $X2=0.5130 $Y2=0.0900
r34 10 21 0.314665 $w=2.27e-07 $l=4.5e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5130 $Y2=0.0900
.ends

.subckt PM_DFFHQNx1_ASAP7_75t_R%SH VSS 11 12 65 68 71 74 28 6 18 14 13 23 25 16
+ 15 17 5 2 22 27 26 20 21 1 24 19
c1 1 VSS 0.000775166f
c2 2 VSS 0.00443737f
c3 5 VSS 0.00500635f
c4 6 VSS 0.0049296f
c5 11 VSS 0.0374582f
c6 12 VSS 0.0801799f
c7 13 VSS 0.00375186f
c8 14 VSS 0.00396971f
c9 15 VSS 0.00862183f
c10 16 VSS 0.00154718f
c11 17 VSS 0.00155981f
c12 18 VSS 0.00220354f
c13 19 VSS 0.000605024f
c14 20 VSS 0.000493736f
c15 21 VSS 0.00100584f
c16 22 VSS 0.00272554f
c17 23 VSS 0.00589929f
c18 24 VSS 0.00230613f
c19 25 VSS 0.000109755f
c20 26 VSS 0.000359629f
c21 27 VSS 0.000317399f
c22 28 VSS 0.00768646f
r1 74 73 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r2 5 73 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6500 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r3 70 5 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6380 $Y=0.0405 $X2=0.6500 $Y2=0.0405
r4 13 70 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0405 $X2=0.6380 $Y2=0.0405
r5 71 13 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.0405 $X2=0.6335 $Y2=0.0405
r6 68 67 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r7 66 67 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7120 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r8 6 66 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7000 $Y=0.2295 $X2=0.7120 $Y2=0.2295
r9 14 6 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.2295 $X2=0.7000 $Y2=0.2295
r10 65 14 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.2295 $X2=0.6875 $Y2=0.2295
r11 5 57 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.0405
+ $X2=0.6480 $Y2=0.0360
r12 2 52 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.9990 $Y=0.1350
+ $X2=0.9990 $Y2=0.1440
r13 12 2 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.9990
+ $Y=0.1350 $X2=0.9990 $Y2=0.1350
r14 6 50 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7020 $Y=0.2295
+ $X2=0.7020 $Y2=0.2330
r15 57 58 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6480
+ $Y=0.0360 $X2=0.6615 $Y2=0.0360
r16 55 58 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0360 $X2=0.6615 $Y2=0.0360
r17 54 55 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6860
+ $Y=0.0360 $X2=0.6750 $Y2=0.0360
r18 15 24 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.7040
+ $Y=0.0360 $X2=0.7290 $Y2=0.0360
r19 15 54 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7040
+ $Y=0.0360 $X2=0.6860 $Y2=0.0360
r20 22 52 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.9990
+ $Y=0.1080 $X2=0.9990 $Y2=0.1440
r21 50 51 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.2330 $X2=0.7155 $Y2=0.2330
r22 23 51 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.2330 $X2=0.7155 $Y2=0.2330
r23 24 43 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.0360 $X2=0.7290 $Y2=0.0630
r24 47 52 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.9990 $Y=0.1530
+ $X2=0.9990 $Y2=0.1440
r25 46 47 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1530 $X2=0.9990 $Y2=0.1530
r26 45 46 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1530 $X2=0.9450 $Y2=0.1530
r27 28 45 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.8795
+ $Y=0.1530 $X2=0.8910 $Y2=0.1530
r28 44 45 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.8910 $Y=0.1485 $X2=0.8910
+ $Y2=0.1530
r29 21 44 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1305 $X2=0.8910 $Y2=0.1485
r30 17 38 6.38362 $w=1.33509e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1975 $X2=0.7290 $Y2=0.1690
r31 17 23 7.09793 $w=1.42676e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1975 $X2=0.7290 $Y2=0.2330
r32 42 43 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.0900 $X2=0.7290 $Y2=0.0630
r33 41 42 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1000 $X2=0.7290 $Y2=0.0900
r34 40 41 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1100 $X2=0.7290 $Y2=0.1000
r35 16 25 4.67854 $w=1.44583e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1360 $X2=0.7290 $Y2=0.1600
r36 16 40 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1360 $X2=0.7290 $Y2=0.1100
r37 27 39 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1575 $X2=0.8910 $Y2=0.1665
r38 27 44 1.50855 $w=1.55e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1575 $X2=0.8910 $Y2=0.1485
r39 27 45 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.8910 $Y=0.1575 $X2=0.8910
+ $Y2=0.1530
r40 25 38 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1600 $X2=0.7290 $Y2=0.1690
r41 37 39 4.19024 $w=1.156e-08 $l=2.54018e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8660 $Y=0.1620 $X2=0.8910 $Y2=0.1665
r42 20 26 1.38478 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8480 $Y=0.1620 $X2=0.8370 $Y2=0.1620
r43 20 37 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8480
+ $Y=0.1620 $X2=0.8660 $Y2=0.1620
r44 36 38 4.4015 $w=1.35e-08 $l=2.78927e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7560 $Y=0.1620 $X2=0.7290 $Y2=0.1690
r45 35 36 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1620 $X2=0.7560 $Y2=0.1620
r46 18 26 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.1620 $X2=0.8370 $Y2=0.1620
r47 18 35 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.1620 $X2=0.7830 $Y2=0.1620
r48 26 34 4.88263 $w=1.47308e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8370 $Y=0.1620 $X2=0.8370 $Y2=0.1360
r49 19 34 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1180 $X2=0.8370 $Y2=0.1360
r50 11 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.8370
+ $Y=0.1350 $X2=0.8370 $Y2=0.1350
r51 1 34 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8370 $Y=0.1350
+ $X2=0.8370 $Y2=0.1360
.ends

.subckt PM_DFFHQNx1_ASAP7_75t_R%PD1 VSS 7 10 5 4 1
c1 1 VSS 0.010626f
c2 4 VSS 0.00319064f
c3 5 VSS 0.00185356f
r1 10 9 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r2 8 9 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r3 5 8 0.123457 $w=8.1e-08 $l=1e-08 $layer=N_src_drn $thickness=1e-09 $X=0.3780
+ $Y=0.0675 $X2=0.3880 $Y2=0.0675
r4 4 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3220 $Y2=0.0675
r5 7 4 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r6 1 5 1e-05
.ends

.subckt PM_DFFHQNx1_ASAP7_75t_R%D VSS 19 3 5 6 7 9 1 4 8
c1 1 VSS 0.010784f
c2 3 VSS 0.0836285f
c3 4 VSS 0.00377208f
c4 5 VSS 0.0034238f
c5 6 VSS 0.00164691f
c6 7 VSS 0.00744815f
c7 8 VSS 0.00111497f
c8 9 VSS 0.00733033f
r1 9 21 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2430 $Y2=0.2140
r2 7 18 5.17411 $w=1.46514e-08 $l=2.72e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0360 $X2=0.2430 $Y2=0.0632
r3 5 8 7.7975 $w=1.41688e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1735 $X2=0.2430 $Y2=0.1350
r4 5 21 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1735 $X2=0.2430 $Y2=0.2140
r5 19 20 2.85657 $w=1.3e-08 $l=1.22e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0820 $X2=0.2430 $Y2=0.0942
r6 19 18 4.37231 $w=1.3e-08 $l=1.88e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0820 $X2=0.2430 $Y2=0.0632
r7 4 8 3.2503 $w=1.53684e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1160 $X2=0.2430 $Y2=0.1350
r8 4 20 5.07188 $w=1.3e-08 $l=2.18e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1160 $X2=0.2430 $Y2=0.0942
r9 16 17 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2715
+ $Y=0.1350 $X2=0.2810 $Y2=0.1350
r10 6 16 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2615
+ $Y=0.1350 $X2=0.2715 $Y2=0.1350
r11 6 8 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2615 $Y=0.1350 $X2=0.2430 $Y2=0.1350
r12 14 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2770 $Y=0.1350
+ $X2=0.2810 $Y2=0.1350
r13 12 14 4.43042 $w=1.53e-08 $l=7.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.2845 $Y=0.1350 $X2=0.2770 $Y2=0.1350
r14 1 11 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.2885
+ $Y=0.1350 $X2=0.2985 $Y2=0.1350
r15 1 12 1.86855 $w=1.78125e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.2885 $Y=0.1350 $X2=0.2845 $Y2=0.1350
r16 3 11 2.53453 $w=1.32811e-07 $l=1.5e-09 $layer=LIG $thickness=5.23243e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2985 $Y2=0.1350
r17 3 12 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2845 $Y2=0.1350
.ends

.subckt PM_DFFHQNx1_ASAP7_75t_R%CLKN VSS 13 14 15 77 79 22 8 26 7 16 17 1 19 21
+ 20 18 28 23 2 24 3
c1 1 VSS 0.00161774f
c2 2 VSS 4.46263e-20
c3 3 VSS 0.000144963f
c4 7 VSS 0.00748533f
c5 8 VSS 0.00761307f
c6 13 VSS 0.0596085f
c7 14 VSS 0.00439492f
c8 15 VSS 0.0045813f
c9 16 VSS 0.00599169f
c10 17 VSS 0.00591866f
c11 18 VSS 0.00529647f
c12 19 VSS 0.00346919f
c13 20 VSS 0.00461664f
c14 21 VSS 0.00450559f
c15 22 VSS 0.000591849f
c16 23 VSS 0.000584764f
c17 24 VSS 0.00139559f
c18 25 VSS 0.0036545f
c19 26 VSS 0.00153761f
c20 27 VSS 0.00379539f
c21 28 VSS 0.0235666f
r1 79 78 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r2 17 78 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r3 77 76 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r4 16 76 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r5 8 74 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0550 $Y2=0.2340
r6 7 71 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0550 $Y2=0.0360
r7 73 74 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.2340 $X2=0.0550 $Y2=0.2340
r8 21 73 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0460 $Y2=0.2340
r9 21 27 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0180 $Y2=0.2340
r10 70 71 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.0360 $X2=0.0550 $Y2=0.0360
r11 20 70 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0460 $Y2=0.0360
r12 20 25 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0180 $Y2=0.0360
r13 27 63 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.2340 $X2=0.0180 $Y2=0.2125
r14 25 61 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.0360 $X2=0.0180 $Y2=0.0575
r15 3 58 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6750 $Y=0.1350
+ $X2=0.6750 $Y2=0.1440
r16 15 3 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6750
+ $Y=0.1350 $X2=0.6750 $Y2=0.1350
r17 2 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
r18 14 2 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r19 62 63 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1820 $X2=0.0180 $Y2=0.2125
r20 19 26 0.998523 $w=1.74118e-08 $l=1.01119e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1630 $X2=0.0165 $Y2=0.1530
r21 19 62 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1630 $X2=0.0180 $Y2=0.1820
r22 60 61 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0880 $X2=0.0180 $Y2=0.0575
r23 18 26 5.19594 $w=1.44151e-08 $l=2.80401e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1250 $X2=0.0165 $Y2=0.1530
r24 18 60 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1250 $X2=0.0180 $Y2=0.0880
r25 24 58 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1135 $X2=0.6750 $Y2=0.1440
r26 23 56 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1530
r27 52 53 1.90199 $w=1.38333e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.0255 $Y=0.1530 $X2=0.0345 $Y2=0.1530
r28 26 52 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0165
+ $Y=0.1530 $X2=0.0255 $Y2=0.1530
r29 50 58 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.6750 $Y=0.1530
+ $X2=0.6750 $Y2=0.1440
r30 49 50 18.3054 $w=1.3e-08 $l=7.85e-08 $layer=M2 $thickness=3.6e-08 $X=0.5965
+ $Y=0.1530 $X2=0.6750 $Y2=0.1530
r31 48 49 29.3819 $w=1.3e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.4705
+ $Y=0.1530 $X2=0.5965 $Y2=0.1530
r32 47 48 15.2739 $w=1.3e-08 $l=6.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1530 $X2=0.4705 $Y2=0.1530
r33 47 56 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4050 $Y=0.1530
+ $X2=0.4050 $Y2=0.1530
r34 46 47 27.8662 $w=1.3e-08 $l=1.195e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.2855 $Y=0.1530 $X2=0.4050 $Y2=0.1530
r35 45 46 27.5164 $w=1.3e-08 $l=1.18e-07 $layer=M2 $thickness=3.6e-08 $X=0.1675
+ $Y=0.1530 $X2=0.2855 $Y2=0.1530
r36 44 45 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M2 $thickness=3.6e-08 $X=0.1510
+ $Y=0.1530 $X2=0.1675 $Y2=0.1530
r37 43 44 13.7582 $w=1.3e-08 $l=5.9e-08 $layer=M2 $thickness=3.6e-08 $X=0.0920
+ $Y=0.1530 $X2=0.1510 $Y2=0.1530
r38 42 43 13.7582 $w=1.3e-08 $l=5.9e-08 $layer=M2 $thickness=3.6e-08 $X=0.0330
+ $Y=0.1530 $X2=0.0920 $Y2=0.1530
r39 42 53 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.0330 $Y=0.1530
+ $X2=0.0345 $Y2=0.1530
r40 28 42 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.0215
+ $Y=0.1530 $X2=0.0330 $Y2=0.1530
r41 39 44 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1510 $Y=0.1440
+ $X2=0.1510 $Y2=0.1530
r42 22 39 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1510
+ $Y=0.1160 $X2=0.1510 $Y2=0.1440
r43 37 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1550 $Y=0.1350
+ $X2=0.1510 $Y2=0.1440
r44 36 37 4.43042 $w=1.53e-08 $l=7.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1475 $Y=0.1350 $X2=0.1550 $Y2=0.1350
r45 34 36 1.86855 $w=1.78125e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1435 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r46 1 34 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.1335
+ $Y=0.1350 $X2=0.1435 $Y2=0.1350
r47 13 1 2.53453 $w=1.32811e-07 $l=1.5e-09 $layer=LIG $thickness=5.23243e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1335 $Y2=0.1350
r48 13 36 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r49 8 17 1e-05
r50 7 16 1e-05
.ends

.subckt PM_DFFHQNx1_ASAP7_75t_R%MH VSS 9 49 53 59 63 10 18 14 12 3 15 4 16 19
+ 17 20 1
c1 1 VSS 0.000361686f
c2 3 VSS 0.00583982f
c3 4 VSS 0.00560408f
c4 9 VSS 0.0363839f
c5 10 VSS 0.00226802f
c6 11 VSS 8.98097e-20
c7 12 VSS 0.00280309f
c8 13 VSS 6.87267e-20
c9 14 VSS 0.00883397f
c10 15 VSS 0.00138593f
c11 16 VSS 0.000721187f
c12 17 VSS 0.000424913f
c13 18 VSS 0.00607497f
c14 19 VSS 1.2099e-20
c15 20 VSS 0.0024007f
r1 63 62 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r2 61 62 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r3 3 61 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3760 $Y=0.2295 $X2=0.3880 $Y2=0.2295
r4 13 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2295 $X2=0.3760 $Y2=0.2295
r5 57 58 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r6 59 57 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.1890 $X2=0.3635 $Y2=0.1890
r7 12 58 0.185185 $w=5.4e-08 $l=1e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r8 12 3 0.518519 $w=3.9e-08 $l=4.05494e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.1890 $X2=0.3760 $Y2=0.2295
r9 3 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2295
+ $X2=0.3780 $Y2=0.2340
r10 53 52 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r11 51 52 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4420 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r12 4 51 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4300 $Y=0.0405 $X2=0.4420 $Y2=0.0405
r13 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0405 $X2=0.4300 $Y2=0.0405
r14 10 4 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0810 $X2=0.4300 $Y2=0.0810
r15 49 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0810 $X2=0.4175 $Y2=0.0810
r16 45 46 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r17 43 46 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r18 42 43 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4160
+ $Y=0.2340 $X2=0.4050 $Y2=0.2340
r19 14 20 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4340
+ $Y=0.2340 $X2=0.4590 $Y2=0.2340
r20 14 42 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4340
+ $Y=0.2340 $X2=0.4160 $Y2=0.2340
r21 4 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0405
+ $X2=0.4320 $Y2=0.0360
r22 20 34 3.01468 $w=1.741e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4590 $Y2=0.2140
r23 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4455 $Y2=0.0360
r24 18 31 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4590 $Y2=0.0630
r25 18 37 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4455 $Y2=0.0360
r26 33 34 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1850 $X2=0.4590 $Y2=0.2140
r27 32 33 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1660 $X2=0.4590 $Y2=0.1850
r28 16 19 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1525 $X2=0.4590 $Y2=0.1310
r29 16 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1525 $X2=0.4590 $Y2=0.1660
r30 30 31 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0900 $X2=0.4590 $Y2=0.0630
r31 29 30 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1025 $X2=0.4590 $Y2=0.0900
r32 15 19 2.78392 $w=1.56471e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1140 $X2=0.4590 $Y2=0.1310
r33 15 29 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1140 $X2=0.4590 $Y2=0.1025
r34 19 28 4.18306 $w=1.49565e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1310 $X2=0.4820 $Y2=0.1310
r35 27 28 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5000
+ $Y=0.1310 $X2=0.4820 $Y2=0.1310
r36 26 27 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1310 $X2=0.5000 $Y2=0.1310
r37 17 25 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1310 $X2=0.5670 $Y2=0.1310
r38 17 26 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1310 $X2=0.5130 $Y2=0.1310
r39 1 22 2.36633 $w=2.3e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.5670
+ $Y=0.1305 $X2=0.5670 $Y2=0.1305
r40 1 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1305
+ $X2=0.5670 $Y2=0.1310
r41 9 22 0.314665 $w=2.27e-07 $l=4.5e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5670 $Y=0.1350 $X2=0.5670 $Y2=0.1305
r42 3 12 1e-05
.ends

.subckt PM_DFFHQNx1_ASAP7_75t_R%CLKB VSS 14 15 16 17 81 83 18 20 26 6 7 23 24 4
+ 25 22 19 1 21 8 2
c1 1 VSS 0.00179857f
c2 2 VSS 0.000806134f
c3 3 VSS 0.000757384f
c4 4 VSS 0.00114283f
c5 6 VSS 0.00886089f
c6 7 VSS 0.00857742f
c7 8 VSS 0.00504955f
c8 14 VSS 0.00605157f
c9 15 VSS 0.00582001f
c10 16 VSS 0.00510313f
c11 17 VSS 0.00593781f
c12 18 VSS 0.00549115f
c13 19 VSS 0.00548471f
c14 20 VSS 0.00411908f
c15 21 VSS 0.003361f
c16 22 VSS 0.00284502f
c17 23 VSS 0.0068745f
c18 24 VSS 0.00608506f
c19 25 VSS 0.00127211f
c20 26 VSS 0.00548518f
r1 19 7 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1600 $Y2=0.2160
r2 83 19 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r3 18 6 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1600 $Y2=0.0540
r4 81 18 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r5 4 79 2.78395 $w=2.4e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08 $X=0.7290
+ $Y=0.1780 $X2=0.7250 $Y2=0.1780
r6 17 4 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.7290 $Y=0.1350 $X2=0.7290 $Y2=0.1780
r7 3 72 10.3807 $w=2.30357e-08 $l=0 $layer=LISD $thickness=3.675e-08 $X=0.6210
+ $Y=0.1780 $X2=0.6210 $Y2=0.1780
r8 16 3 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.6210 $Y=0.1350 $X2=0.6210 $Y2=0.1780
r9 2 65 2.78395 $w=2.4e-08 $l=5e-09 $layer=LIG $thickness=4.8e-08 $X=0.4590
+ $Y=0.1780 $X2=0.4640 $Y2=0.1780
r10 15 2 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4590 $Y2=0.1780
r11 7 57 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1655 $Y2=0.2340
r12 6 53 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1655 $Y2=0.0360
r13 78 79 4.8113 $w=2.22e-08 $l=1.5e-09 $layer=LISD $thickness=2.7e-08
+ $X=0.7235 $Y=0.1780 $X2=0.7250 $Y2=0.1780
r14 77 78 10.8887 $w=2.22e-08 $l=2.15e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7020 $Y=0.1780 $X2=0.7235 $Y2=0.1780
r15 76 77 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6885 $Y=0.1780 $X2=0.7020 $Y2=0.1780
r16 75 76 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6750 $Y=0.1780 $X2=0.6885 $Y2=0.1780
r17 74 75 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6615 $Y=0.1780 $X2=0.6750 $Y2=0.1780
r18 73 74 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6480 $Y=0.1780 $X2=0.6615 $Y2=0.1780
r19 72 73 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6210 $Y=0.1780 $X2=0.6480 $Y2=0.1780
r20 71 72 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5940 $Y=0.1780 $X2=0.6210 $Y2=0.1780
r21 70 71 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5805 $Y=0.1780 $X2=0.5940 $Y2=0.1780
r22 69 70 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5670 $Y=0.1780 $X2=0.5805 $Y2=0.1780
r23 68 69 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5535 $Y=0.1780 $X2=0.5670 $Y2=0.1780
r24 67 68 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5400 $Y=0.1780 $X2=0.5535 $Y2=0.1780
r25 66 67 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5265 $Y=0.1780 $X2=0.5400 $Y2=0.1780
r26 64 65 10.3823 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4775 $Y=0.1780 $X2=0.4640 $Y2=0.1780
r27 63 64 11.142 $w=2.22e-08 $l=2.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4995 $Y=0.1780 $X2=0.4775 $Y2=0.1780
r28 62 66 1.51936 $w=2.22e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.5235
+ $Y=0.1780 $X2=0.5265 $Y2=0.1780
r29 61 62 5.31775 $w=2.22e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5130 $Y=0.1780 $X2=0.5235 $Y2=0.1780
r30 8 61 5.31775 $w=2.22e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5025 $Y=0.1780 $X2=0.5130 $Y2=0.1780
r31 8 63 1.51936 $w=2.22e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.5025
+ $Y=0.1780 $X2=0.4995 $Y2=0.1780
r32 57 58 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1655
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r33 24 50 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2340 $X2=0.1890 $Y2=0.2125
r34 24 58 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2340 $X2=0.1755 $Y2=0.2340
r35 53 54 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1655
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r36 23 49 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1890 $Y2=0.0575
r37 23 54 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1755 $Y2=0.0360
r38 51 61 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5130 $Y=0.1845
+ $X2=0.5130 $Y2=0.1780
r39 22 51 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1680 $X2=0.5130 $Y2=0.1845
r40 48 49 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0880 $X2=0.1890 $Y2=0.0575
r41 47 48 11.3097 $w=1.3e-08 $l=4.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1365 $X2=0.1890 $Y2=0.0880
r42 46 50 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1990 $X2=0.1890 $Y2=0.2125
r43 45 46 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1890 $X2=0.1890 $Y2=0.1990
r44 20 45 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1735 $X2=0.1890 $Y2=0.1890
r45 20 47 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1735 $X2=0.1890 $Y2=0.1365
r46 43 51 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.5130 $Y=0.1890
+ $X2=0.5130 $Y2=0.1845
r47 42 43 22.0364 $w=1.3e-08 $l=9.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.4185
+ $Y=0.1890 $X2=0.5130 $Y2=0.1890
r48 41 42 22.0364 $w=1.3e-08 $l=9.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1890 $X2=0.4185 $Y2=0.1890
r49 40 41 15.7403 $w=1.3e-08 $l=6.75e-08 $layer=M2 $thickness=3.6e-08 $X=0.2565
+ $Y=0.1890 $X2=0.3240 $Y2=0.1890
r50 39 40 15.7403 $w=1.3e-08 $l=6.75e-08 $layer=M2 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1890 $X2=0.2565 $Y2=0.1890
r51 39 45 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1890 $Y=0.1890
+ $X2=0.1890 $Y2=0.1890
r52 26 39 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.1775
+ $Y=0.1890 $X2=0.1890 $Y2=0.1890
r53 37 41 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.3240 $Y=0.1890
+ $X2=0.3240 $Y2=0.1890
r54 36 37 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1735 $X2=0.3240 $Y2=0.1890
r55 21 34 3.60008 $w=1.51951e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3240 $Y=0.1555 $X2=0.3240 $Y2=0.1350
r56 21 36 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1555 $X2=0.3240 $Y2=0.1735
r57 25 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r58 25 34 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3375 $Y=0.1350 $X2=0.3240 $Y2=0.1350
r59 14 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r60 1 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
.ends


*
.SUBCKT DFFHQNx1_ASAP7_75t_R VSS VDD CLK D QN
*
* VSS VSS
* VDD VDD
* CLK CLK
* D D
* QN QN
*
*

MM20 N_MM20_d N_MM20_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM23 N_MM23_d N_MM22_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM10_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM6 N_MM6_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM12 N_MM12_d N_MM12_g N_MM12_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM17 N_MM17_d N_MM13_g N_MM17_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM16 N_MM16_d N_MM19_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM14 N_MM14_d N_MM14_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM24 N_MM24_d N_MM24_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM21 N_MM21_d N_MM20_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM22 N_MM22_d N_MM22_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM13 N_MM13_d N_MM13_g N_MM13_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM18 N_MM18_d N_MM18_g N_MM18_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM19 N_MM19_d N_MM19_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM15 N_MM15_d N_MM14_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM25 N_MM25_d N_MM24_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "DFFHQNx1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "DFFHQNx1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_DFFHQNx1_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_DFFHQNx1_ASAP7_75t_R%noxref_18
cc_1 N_noxref_18_1 N_MM20_g 0.00368344f
cc_2 N_noxref_18_1 N_CLKN_19 6.2419e-20
cc_3 N_noxref_18_1 N_CLKN_18 0.000313322f
cc_4 N_noxref_18_1 N_CLKN_7 0.000503374f
cc_5 N_noxref_18_1 N_CLKN_16 0.027831f
x_PM_DFFHQNx1_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_DFFHQNx1_ASAP7_75t_R%noxref_19
cc_6 N_noxref_19_1 N_MM20_g 0.00367249f
cc_7 N_noxref_19_1 N_CLKN_26 8.87656e-20
cc_8 N_noxref_19_1 N_CLKN_18 0.0001526f
cc_9 N_noxref_19_1 N_CLKN_19 0.000196767f
cc_10 N_noxref_19_1 N_CLKN_8 0.000505002f
cc_11 N_noxref_19_1 N_CLKN_17 0.0278538f
cc_12 N_noxref_19_1 N_noxref_18_1 0.00204872f
x_PM_DFFHQNx1_ASAP7_75t_R%noxref_29 VSS N_noxref_29_1
+ PM_DFFHQNx1_ASAP7_75t_R%noxref_29
cc_13 N_noxref_29_1 N_MM24_g 0.00148788f
cc_14 N_noxref_29_1 N_QN_8 0.0385712f
cc_15 N_noxref_29_1 N_noxref_28_1 0.00177171f
x_PM_DFFHQNx1_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_DFFHQNx1_ASAP7_75t_R%noxref_24
cc_16 N_noxref_24_1 N_SS_10 0.017019f
cc_17 N_noxref_24_1 N_MM14_g 0.00610649f
x_PM_DFFHQNx1_ASAP7_75t_R%noxref_28 VSS N_noxref_28_1
+ PM_DFFHQNx1_ASAP7_75t_R%noxref_28
cc_18 N_noxref_28_1 N_MM24_g 0.00148998f
cc_19 N_noxref_28_1 N_QN_7 0.0383584f
x_PM_DFFHQNx1_ASAP7_75t_R%noxref_26 VSS N_noxref_26_1
+ PM_DFFHQNx1_ASAP7_75t_R%noxref_26
cc_20 N_noxref_26_1 N_SS_10 0.00063801f
cc_21 N_noxref_26_1 N_MM24_g 0.00169018f
cc_22 N_noxref_26_1 N_noxref_24_1 0.00776243f
cc_23 N_noxref_26_1 N_noxref_25_1 0.000480418f
x_PM_DFFHQNx1_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_DFFHQNx1_ASAP7_75t_R%noxref_25
cc_24 N_noxref_25_1 N_SS_11 0.0169303f
cc_25 N_noxref_25_1 N_SH_1 0.000200845f
cc_26 N_noxref_25_1 N_MM14_g 0.00600389f
cc_27 N_noxref_25_1 N_noxref_24_1 0.00152869f
x_PM_DFFHQNx1_ASAP7_75t_R%noxref_27 VSS N_noxref_27_1
+ PM_DFFHQNx1_ASAP7_75t_R%noxref_27
cc_28 N_noxref_27_1 N_SS_11 0.000629057f
cc_29 N_noxref_27_1 N_MM24_g 0.0017122f
cc_30 N_noxref_27_1 N_noxref_24_1 0.000482892f
cc_31 N_noxref_27_1 N_noxref_25_1 0.00775912f
cc_32 N_noxref_27_1 N_noxref_26_1 0.00124004f
x_PM_DFFHQNx1_ASAP7_75t_R%QN VSS QN N_MM24_d N_MM25_d N_QN_2 N_QN_7 N_QN_9
+ N_QN_1 N_QN_8 PM_DFFHQNx1_ASAP7_75t_R%QN
cc_33 N_QN_2 N_SS_17 0.000428839f
cc_34 N_QN_2 N_SS_15 0.00179808f
cc_35 N_QN_7 N_SH_22 0.00111255f
cc_36 N_QN_9 N_SH_28 0.000838168f
cc_37 N_QN_2 N_SH_2 0.000895953f
cc_38 N_QN_2 N_MM24_g 0.00117365f
cc_39 N_QN_1 N_MM24_g 0.00124412f
cc_40 N_QN_8 N_SH_2 0.00173727f
cc_41 N_QN_9 N_SH_22 0.00547407f
cc_42 N_QN_8 N_MM24_g 0.0154663f
cc_43 N_QN_7 N_MM24_g 0.0543398f
x_PM_DFFHQNx1_ASAP7_75t_R%PD3 VSS N_MM9_s N_MM8_d N_PD3_1
+ PM_DFFHQNx1_ASAP7_75t_R%PD3
cc_44 N_PD3_1 N_MM9_g 0.00773025f
cc_45 N_PD3_1 N_MM11_g 0.00773412f
x_PM_DFFHQNx1_ASAP7_75t_R%PD4 VSS N_MM18_s N_MM19_d N_PD4_1
+ PM_DFFHQNx1_ASAP7_75t_R%PD4
cc_46 N_PD4_1 N_MM18_g 0.00773069f
cc_47 N_PD4_1 N_MM19_g 0.00776505f
x_PM_DFFHQNx1_ASAP7_75t_R%PU1 VSS N_MM3_d N_MM1_s N_PU1_1
+ PM_DFFHQNx1_ASAP7_75t_R%PU1
cc_48 N_PU1_1 N_MM3_g 0.0171024f
cc_49 N_PU1_1 N_MM1_g 0.0169758f
x_PM_DFFHQNx1_ASAP7_75t_R%PD2 VSS N_MM10_s N_MM11_d N_PD2_4 N_PD2_5 N_PD2_1
+ PM_DFFHQNx1_ASAP7_75t_R%PD2
cc_50 N_PD2_4 N_MM10_g 0.0150486f
cc_51 N_PD2_5 N_CLKB_8 0.00146961f
cc_52 N_PD2_1 N_CLKB_2 0.000539914f
cc_53 N_PD2_1 N_MM9_g 0.0020622f
cc_54 N_PD2_4 N_MM9_g 0.00714095f
cc_55 N_PD2_5 N_MM9_g 0.0240567f
cc_56 N_PD2_5 N_MM11_g 0.014603f
cc_57 N_PD2_1 N_MH_14 0.00043568f
cc_58 N_PD2_4 N_MH_3 0.000614553f
cc_59 N_PD2_1 N_MH_20 0.00320688f
x_PM_DFFHQNx1_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_DFFHQNx1_ASAP7_75t_R%noxref_20
cc_60 N_noxref_20_1 N_CLKN_1 0.000398066f
cc_61 N_noxref_20_1 N_MM22_g 0.00343386f
cc_62 N_noxref_20_1 N_CLKB_6 0.000423111f
cc_63 N_noxref_20_1 N_CLKB_18 0.0270305f
x_PM_DFFHQNx1_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_DFFHQNx1_ASAP7_75t_R%noxref_22
cc_64 N_noxref_22_1 N_MM3_g 0.00183864f
cc_65 N_noxref_22_1 N_CLKB_6 0.000104326f
cc_66 N_noxref_22_1 N_CLKB_18 0.000553087f
cc_67 N_noxref_22_1 N_noxref_20_1 0.00768743f
cc_68 N_noxref_22_1 N_noxref_21_1 0.000463733f
x_PM_DFFHQNx1_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_DFFHQNx1_ASAP7_75t_R%noxref_21
cc_69 N_noxref_21_1 N_CLKN_1 0.000396541f
cc_70 N_noxref_21_1 N_MM22_g 0.00344681f
cc_71 N_noxref_21_1 N_CLKB_7 0.000426471f
cc_72 N_noxref_21_1 N_CLKB_19 0.0270305f
cc_73 N_noxref_21_1 N_noxref_20_1 0.00141787f
x_PM_DFFHQNx1_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_DFFHQNx1_ASAP7_75t_R%noxref_23
cc_74 N_noxref_23_1 N_MM3_g 0.0018533f
cc_75 N_noxref_23_1 N_CLKB_7 0.000100589f
cc_76 N_noxref_23_1 N_CLKB_19 0.000556467f
cc_77 N_noxref_23_1 N_noxref_20_1 0.000463245f
cc_78 N_noxref_23_1 N_noxref_21_1 0.00768972f
cc_79 N_noxref_23_1 N_noxref_22_1 0.00122256f
x_PM_DFFHQNx1_ASAP7_75t_R%SS VSS N_MM19_g N_MM14_d N_MM15_d N_SS_12 N_SS_10
+ N_SS_11 N_SS_15 N_SS_4 N_SS_3 N_SS_14 N_SS_1 N_SS_16 N_SS_13 N_SS_17
+ PM_DFFHQNx1_ASAP7_75t_R%SS
cc_80 N_MM19_g N_CLKB_8 0.000215376f
cc_81 N_MM19_g N_CLKB_4 0.000537906f
cc_82 N_MM19_g N_MM18_g 0.0135231f
x_PM_DFFHQNx1_ASAP7_75t_R%PD5 VSS N_MM17_s N_MM16_d N_PD5_4 N_PD5_1 N_PD5_5
+ PM_DFFHQNx1_ASAP7_75t_R%PD5
cc_83 N_PD5_4 N_MM13_g 0.0152724f
cc_84 N_PD5_1 N_MM18_g 0.000759519f
cc_85 N_PD5_4 N_MM18_g 0.00695235f
cc_86 N_PD5_5 N_MM18_g 0.023986f
cc_87 N_PD5_1 N_MM19_g 0.000916096f
cc_88 N_PD5_5 N_MM19_g 0.0155328f
cc_89 N_PD5_1 N_SH_13 0.000516336f
cc_90 N_PD5_1 N_SH_15 0.000437004f
cc_91 N_PD5_1 N_SH_16 0.000599659f
cc_92 N_PD5_4 N_SH_5 0.000664456f
cc_93 N_PD5_1 N_SH_24 0.00238016f
x_PM_DFFHQNx1_ASAP7_75t_R%CLK VSS CLK N_MM20_g N_CLK_8 N_CLK_5 N_CLK_1 N_CLK_6
+ N_CLK_7 N_CLK_4 PM_DFFHQNx1_ASAP7_75t_R%CLK
x_PM_DFFHQNx1_ASAP7_75t_R%MS VSS N_MM11_g N_MM6_d N_MM12_d N_MM7_d N_MM13_d
+ N_MS_13 N_MS_17 N_MS_18 N_MS_14 N_MS_3 N_MS_15 N_MS_12 N_MS_1 N_MS_11 N_MS_4
+ N_MS_16 PM_DFFHQNx1_ASAP7_75t_R%MS
cc_94 N_MS_13 N_MM10_g 0.000130138f
cc_95 N_MS_13 N_CLKN_24 0.00032756f
cc_96 N_MS_13 N_CLKN_28 0.00022929f
cc_97 N_MS_13 N_CLKN_3 0.000229581f
cc_98 N_MS_17 N_CLKN_24 0.00452728f
cc_99 N_MS_17 N_CLKN_3 0.000282384f
cc_100 N_MS_18 N_CLKN_24 0.000632715f
cc_101 N_MS_14 N_CLKN_28 0.00276276f
cc_102 N_MS_13 N_MM13_g 0.0153408f
cc_103 N_MS_3 N_CLKB_8 0.00055579f
cc_104 N_MS_3 N_CLKB_2 0.000123737f
cc_105 N_MS_3 N_CLKB_22 0.000154806f
cc_106 N_MS_3 N_MM9_g 0.000165533f
cc_107 N_MS_3 N_CLKB_26 0.000172145f
cc_108 N_MS_15 N_CLKB_22 0.000290783f
cc_109 N_MS_12 N_MM12_g 0.0078041f
cc_110 N_MS_13 N_MM12_g 0.00777346f
cc_111 N_MS_15 N_CLKB_8 0.000383383f
cc_112 N_MS_1 N_MM9_g 0.000560232f
cc_113 N_MS_17 N_CLKB_8 0.00157515f
cc_114 N_MS_11 N_MM12_g 0.00651789f
cc_115 N_MS_4 N_MM12_g 0.00255242f
cc_116 N_MS_4 N_CLKB_8 0.00635858f
cc_117 N_MM11_g N_MM9_g 0.0142056f
cc_118 N_MS_3 N_MM12_g 0.0259332f
x_PM_DFFHQNx1_ASAP7_75t_R%SH VSS N_MM14_g N_MM24_g N_MM13_s N_MM18_d N_MM12_s
+ N_MM17_d N_SH_28 N_SH_6 N_SH_18 N_SH_14 N_SH_13 N_SH_23 N_SH_25 N_SH_16
+ N_SH_15 N_SH_17 N_SH_5 N_SH_2 N_SH_22 N_SH_27 N_SH_26 N_SH_20 N_SH_21 N_SH_1
+ N_SH_24 N_SH_19 PM_DFFHQNx1_ASAP7_75t_R%SH
cc_119 N_SH_28 N_CLKN_28 0.000146396f
cc_120 N_SH_6 N_MM13_g 0.000163831f
cc_121 N_SH_18 N_CLKN_24 0.000215659f
cc_122 N_SH_14 N_MM13_g 0.00675259f
cc_123 N_SH_13 N_MM13_g 0.0067885f
cc_124 N_SH_23 N_CLKN_24 0.000362f
cc_125 N_SH_25 N_CLKN_24 0.000937135f
cc_126 N_SH_16 N_CLKN_3 0.000445115f
cc_127 N_SH_15 N_CLKN_24 0.000508874f
cc_128 N_SH_17 N_CLKN_24 0.00052299f
cc_129 N_SH_5 N_CLKN_3 0.000536728f
cc_130 N_SH_15 N_CLKN_28 0.00110287f
cc_131 N_SH_16 N_CLKN_24 0.00388659f
cc_132 N_SH_5 N_MM13_g 0.0184186f
cc_133 N_SH_14 N_CLKB_26 8.72929e-20
cc_134 N_SH_23 N_CLKB_8 0.000188313f
cc_135 N_SH_25 N_CLKB_8 0.000201135f
cc_136 N_SH_13 N_MM12_g 0.00677653f
cc_137 N_SH_6 N_CLKB_8 0.000297547f
cc_138 N_SH_18 N_CLKB_4 0.000403842f
cc_139 N_SH_16 N_CLKB_8 0.000420064f
cc_140 N_SH_17 N_CLKB_8 0.000613358f
cc_141 N_SH_14 N_CLKB_4 0.000928311f
cc_142 N_SH_6 N_MM18_g 0.000989101f
cc_143 N_SH_14 N_CLKB_8 0.00230339f
cc_144 N_SH_5 N_MM12_g 0.0095145f
cc_145 N_SH_14 N_MM18_g 0.0162713f
cc_146 N_SH_16 N_MS_3 0.000112263f
cc_147 N_SH_23 N_MS_3 0.00013281f
cc_148 N_SH_6 N_MS_3 0.000211236f
cc_149 N_SH_14 N_MS_3 0.000438565f
cc_150 N_SH_13 N_MS_3 0.000463915f
cc_151 N_SH_23 N_MS_4 0.000297153f
cc_152 N_SH_6 N_MS_4 0.000418085f
cc_153 N_SH_15 N_MS_16 0.000459173f
cc_154 N_SH_14 N_MS_4 0.000582695f
cc_155 N_SH_23 N_MS_17 0.000613579f
cc_156 N_SH_15 N_MS_18 0.00163754f
cc_157 N_SH_5 N_MS_3 0.00380041f
cc_158 N_SH_2 N_MM19_g 0.000136132f
cc_159 N_SH_17 N_MM19_g 0.000140348f
cc_160 N_SH_22 N_MM19_g 0.00019066f
cc_161 N_SH_27 N_MM19_g 0.000199208f
cc_162 N_SH_26 N_SS_12 0.000215496f
cc_163 N_MM14_g N_SS_10 0.00686392f
cc_164 N_MM14_g N_SS_11 0.00683173f
cc_165 N_SH_22 N_SS_15 0.00713324f
cc_166 N_SH_2 N_SS_15 0.00028578f
cc_167 N_SH_20 N_SS_4 0.000330635f
cc_168 N_SH_21 N_SS_15 0.00181662f
cc_169 N_MM14_g N_SS_3 0.000397637f
cc_170 N_MM14_g N_SS_4 0.000516529f
cc_171 N_SH_20 N_SS_14 0.000650473f
cc_172 N_SH_1 N_SS_1 0.000686419f
cc_173 N_SH_24 N_SS_16 0.000794357f
cc_174 N_SH_16 N_SS_1 0.000849146f
cc_175 N_SH_27 N_SS_15 0.000900288f
cc_176 N_SH_19 N_SS_12 0.000940836f
cc_177 N_SH_21 N_SS_13 0.00106197f
cc_178 N_MM14_g N_SS_1 0.00113556f
cc_179 N_SH_27 N_SS_14 0.00125914f
cc_180 N_SH_1 N_MM19_g 0.00129566f
cc_181 N_SH_18 N_SS_12 0.00159478f
cc_182 N_SH_28 N_SS_15 0.00187091f
cc_183 N_SH_16 N_SS_12 0.00473107f
cc_184 N_MM14_g N_MM19_g 0.0294458f
x_PM_DFFHQNx1_ASAP7_75t_R%PD1 VSS N_MM5_d N_MM4_s N_PD1_5 N_PD1_4 N_PD1_1
+ PM_DFFHQNx1_ASAP7_75t_R%PD1
cc_185 N_PD1_5 N_CLKN_2 0.000858338f
cc_186 N_PD1_5 N_CLKN_23 0.00031664f
cc_187 N_PD1_5 N_MM10_g 0.0343258f
cc_188 N_PD1_4 N_MM3_g 0.0359349f
cc_189 N_PD1_5 N_CLKB_25 0.000412994f
cc_190 N_PD1_5 N_CLKB_1 0.00234462f
cc_191 N_PD1_5 N_MM1_g 0.0735596f
cc_192 N_PD1_1 N_MH_4 0.00122236f
cc_193 N_PD1_1 N_MH_10 0.00350006f
x_PM_DFFHQNx1_ASAP7_75t_R%D VSS D N_MM3_g N_D_5 N_D_6 N_D_7 N_D_9 N_D_1 N_D_4
+ N_D_8 PM_DFFHQNx1_ASAP7_75t_R%D
cc_194 N_D_5 N_CLKN_22 0.000146036f
cc_195 N_D_5 N_CLKN_23 7.47542e-20
cc_196 N_D_5 N_CLKN_1 0.000102901f
cc_197 N_D_6 N_CLKN_28 0.000657125f
cc_198 N_D_5 N_CLKN_28 0.00330948f
x_PM_DFFHQNx1_ASAP7_75t_R%CLKN VSS N_MM22_g N_MM10_g N_MM13_g N_MM20_d N_MM21_d
+ N_CLKN_22 N_CLKN_8 N_CLKN_26 N_CLKN_7 N_CLKN_16 N_CLKN_17 N_CLKN_1 N_CLKN_19
+ N_CLKN_21 N_CLKN_20 N_CLKN_18 N_CLKN_28 N_CLKN_23 N_CLKN_2 N_CLKN_24 N_CLKN_3
+ PM_DFFHQNx1_ASAP7_75t_R%CLKN
cc_199 N_CLKN_22 N_MM20_g 0.000243475f
cc_200 N_CLKN_8 N_MM20_g 0.00112888f
cc_201 N_CLKN_26 N_MM20_g 0.000258164f
cc_202 N_CLKN_7 N_MM20_g 0.0011647f
cc_203 N_CLKN_16 N_MM20_g 0.0112193f
cc_204 N_CLKN_17 N_MM20_g 0.0113277f
cc_205 N_CLKN_1 N_CLK_8 0.000441582f
cc_206 N_CLKN_19 N_CLK_8 0.000504395f
cc_207 N_CLKN_21 N_CLK_8 0.000765329f
cc_208 N_CLKN_20 N_CLK_5 0.000800078f
cc_209 N_CLKN_26 N_CLK_1 0.000803931f
cc_210 N_CLKN_21 N_CLK_6 0.000842599f
cc_211 N_CLKN_22 N_CLK_7 0.001063f
cc_212 N_CLKN_18 N_CLK_7 0.00116006f
cc_213 N_CLKN_26 N_CLK_8 0.00178252f
cc_214 N_CLKN_28 N_CLK_8 0.0018027f
cc_215 N_CLKN_1 N_CLK_1 0.00248534f
cc_216 N_CLKN_20 N_CLK_7 0.00268142f
cc_217 N_CLKN_22 N_CLK_8 0.00324624f
cc_218 N_CLKN_26 N_CLK_4 0.00343261f
cc_219 N_MM22_g N_MM20_g 0.0350526f
x_PM_DFFHQNx1_ASAP7_75t_R%MH VSS N_MM7_g N_MM4_d N_MM9_d N_MM1_d N_MM10_d
+ N_MH_10 N_MH_18 N_MH_14 N_MH_12 N_MH_3 N_MH_15 N_MH_4 N_MH_16 N_MH_19 N_MH_17
+ N_MH_20 N_MH_1 PM_DFFHQNx1_ASAP7_75t_R%MH
cc_220 N_MH_10 N_CLKN_3 0.000103908f
cc_221 N_MH_10 N_CLKN_28 0.000110957f
cc_222 N_MH_10 N_MM13_g 0.000188912f
cc_223 N_MH_10 N_CLKN_23 0.000326487f
cc_224 N_MH_18 N_CLKN_23 0.000369631f
cc_225 N_MH_14 N_CLKN_23 0.000395921f
cc_226 N_MH_12 N_MM10_g 0.0164209f
cc_227 N_MH_3 N_CLKN_2 0.000773564f
cc_228 N_MH_15 N_CLKN_23 0.00110431f
cc_229 N_MH_4 N_MM10_g 0.00111931f
cc_230 N_MH_3 N_MM10_g 0.00123205f
cc_231 N_MH_16 N_CLKN_23 0.00124312f
cc_232 N_MH_10 N_CLKN_2 0.00164702f
cc_233 N_MH_19 N_CLKN_23 0.00296551f
cc_234 N_MH_17 N_CLKN_28 0.00352163f
cc_235 N_MH_10 N_MM10_g 0.0529625f
cc_236 N_MH_10 N_CLKB_22 0.000365904f
cc_237 N_MH_10 N_MM1_g 0.000402116f
cc_238 N_MH_10 N_CLKB_21 0.000176925f
cc_239 N_MH_10 N_CLKB_25 0.000272549f
cc_240 N_MH_20 N_CLKB_22 0.000316083f
cc_241 N_MH_16 N_CLKB_22 0.00266629f
cc_242 N_MH_3 N_CLKB_1 0.000337909f
cc_243 N_MH_17 N_CLKB_8 0.000557181f
cc_244 N_MH_4 N_MM9_g 0.000623346f
cc_245 N_MH_3 N_CLKB_21 0.000652262f
cc_246 N_MH_1 N_CLKB_8 0.0022732f
cc_247 N_MH_16 N_CLKB_2 0.000779051f
cc_248 N_MH_12 N_CLKB_1 0.000794379f
cc_249 N_MH_3 N_MM1_g 0.00175407f
cc_250 N_MH_14 N_CLKB_26 0.00280082f
cc_251 N_MH_17 N_CLKB_22 0.00357875f
cc_252 N_MM7_g N_CLKB_8 0.00464711f
cc_253 N_MH_12 N_MM1_g 0.0336879f
cc_254 N_MM7_g N_MM12_g 0.0127392f
cc_255 N_MH_10 N_MM9_g 0.0363982f
cc_256 N_MH_17 N_MM11_g 0.000358784f
cc_257 N_MH_4 N_MS_1 0.000395618f
cc_258 N_MH_17 N_MS_1 0.000829497f
cc_259 N_MM7_g N_MS_3 0.000906387f
cc_260 N_MH_1 N_MS_14 0.000924544f
cc_261 N_MH_17 N_MS_17 0.00101601f
cc_262 N_MH_1 N_MM11_g 0.00114137f
cc_263 N_MM7_g N_MS_1 0.00116068f
cc_264 N_MH_15 N_MS_14 0.00124156f
cc_265 N_MM7_g N_MS_12 0.00639117f
cc_266 N_MM7_g N_MS_11 0.00640924f
cc_267 N_MH_17 N_MS_14 0.00746951f
cc_268 N_MM7_g N_MM11_g 0.0293597f
x_PM_DFFHQNx1_ASAP7_75t_R%CLKB VSS N_MM1_g N_MM9_g N_MM12_g N_MM18_g N_MM23_d
+ N_MM22_d N_CLKB_18 N_CLKB_20 N_CLKB_26 N_CLKB_6 N_CLKB_7 N_CLKB_23 N_CLKB_24
+ N_CLKB_4 N_CLKB_25 N_CLKB_22 N_CLKB_19 N_CLKB_1 N_CLKB_21 N_CLKB_8 N_CLKB_2
+ PM_DFFHQNx1_ASAP7_75t_R%CLKB
cc_269 N_CLKB_18 N_CLK_6 8.57854e-20
cc_270 N_CLKB_20 N_CLK_6 9.12674e-20
cc_271 N_CLKB_26 N_CLK_6 0.000123345f
cc_272 N_CLKB_6 N_CLK_6 0.000361693f
cc_273 N_CLKB_7 N_CLK_6 0.000387298f
cc_274 N_CLKB_23 N_CLK_7 0.000500038f
cc_275 N_CLKB_20 N_CLK_8 0.000514705f
cc_276 N_CLKB_23 N_CLK_5 0.00120151f
cc_277 N_CLKB_24 N_CLK_6 0.00199622f
cc_278 N_CLKB_6 N_MM22_g 0.000721222f
cc_279 N_CLKB_7 N_MM22_g 0.000747071f
cc_280 N_CLKB_4 N_MM13_g 0.000222558f
cc_281 N_CLKB_25 N_CLKN_28 0.000285919f
cc_282 N_CLKB_22 N_CLKN_28 0.000669652f
cc_283 N_CLKB_24 N_CLKN_22 0.000310766f
cc_284 N_CLKB_19 N_MM22_g 0.0110945f
cc_285 N_CLKB_23 N_CLKN_22 0.000357496f
cc_286 N_CLKB_1 N_CLKN_2 0.00169517f
cc_287 N_CLKB_21 N_CLKN_28 0.00104596f
cc_288 N_CLKB_20 N_CLKN_22 0.00766508f
cc_289 N_CLKB_20 N_CLKN_28 0.000519084f
cc_290 N_CLKB_8 N_CLKN_24 0.000534456f
cc_291 N_CLKB_25 N_CLKN_2 0.000549016f
cc_292 N_CLKB_2 N_MM10_g 0.000589093f
cc_293 N_CLKB_26 N_CLKN_23 0.000616959f
cc_294 N_CLKB_8 N_CLKN_3 0.00279616f
cc_295 N_CLKB_20 N_CLKN_1 0.000691464f
cc_296 N_CLKB_19 N_CLKN_1 0.00121517f
cc_297 N_MM1_g N_MM10_g 0.00164352f
cc_298 N_CLKB_25 N_CLKN_23 0.00263609f
cc_299 N_CLKB_8 N_MM13_g 0.00423843f
cc_300 N_MM12_g N_MM13_g 0.0057225f
cc_301 N_MM9_g N_MM10_g 0.00910615f
cc_302 N_MM18_g N_MM13_g 0.0184454f
cc_303 N_CLKB_26 N_CLKN_28 0.0306005f
cc_304 N_CLKB_18 N_MM22_g 0.0389029f
cc_305 N_CLKB_6 N_MM3_g 0.00011685f
cc_306 N_CLKB_21 N_MM3_g 0.000132909f
cc_307 N_CLKB_20 N_MM3_g 0.000186961f
cc_308 N_CLKB_1 N_MM3_g 0.000265584f
cc_309 N_CLKB_25 N_MM3_g 0.000617636f
cc_310 N_CLKB_23 N_D_7 0.000854403f
cc_311 N_CLKB_26 N_D_6 0.00108917f
cc_312 N_CLKB_21 N_D_6 0.0011142f
cc_313 N_CLKB_24 N_D_9 0.00121817f
cc_314 N_CLKB_1 N_D_1 0.00161854f
cc_315 N_CLKB_20 N_D_4 0.00180992f
cc_316 N_CLKB_25 N_D_6 0.00203563f
cc_317 N_CLKB_20 N_D_5 0.00266241f
cc_318 N_CLKB_20 N_D_8 0.00411765f
cc_319 N_MM1_g N_MM3_g 0.00527925f
*END of DFFHQNx1_ASAP7_75t_R.pxi
.ENDS
** Design:	DFFHQNx2_ASAP7_75t_R
* Created:	"Fri Aug 17 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "DFFHQNx2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "DFFHQNx2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_DFFHQNx2_ASAP7_75t_R%PD3 VSS 2 4 1
c1 1 VSS 0.000972282f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0405 $X2=0.4905 $Y2=0.0405
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0405 $X2=0.4735 $Y2=0.0405
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4735 $Y=0.0405 $X2=0.4905 $Y2=0.0405
.ends

.subckt PM_DFFHQNx2_ASAP7_75t_R%PU1 VSS 2 4 1
c1 1 VSS 0.000984732f
r1 4 3 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3365 $Y2=0.2025
r2 2 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3195 $Y2=0.2025
r3 1 3 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3195 $Y=0.2025 $X2=0.3365 $Y2=0.2025
.ends

.subckt PM_DFFHQNx2_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.0415702f
.ends

.subckt PM_DFFHQNx2_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.0415594f
.ends

.subckt PM_DFFHQNx2_ASAP7_75t_R%PD4 VSS 2 4 1
c1 1 VSS 0.00094577f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.2295 $X2=0.7605 $Y2=0.2295
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.2295 $X2=0.7435 $Y2=0.2295
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7435 $Y=0.2295 $X2=0.7605 $Y2=0.2295
.ends

.subckt PM_DFFHQNx2_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.00426225f
.ends

.subckt PM_DFFHQNx2_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.00486995f
.ends

.subckt PM_DFFHQNx2_ASAP7_75t_R%D VSS 19 3 5 6 7 9 1 4 8
c1 1 VSS 0.0107786f
c2 3 VSS 0.083629f
c3 4 VSS 0.0037761f
c4 5 VSS 0.00342415f
c5 6 VSS 0.00164726f
c6 7 VSS 0.00744929f
c7 8 VSS 0.00111531f
c8 9 VSS 0.00732428f
r1 9 21 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2430 $Y2=0.2140
r2 7 18 5.17411 $w=1.46514e-08 $l=2.72e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0360 $X2=0.2430 $Y2=0.0632
r3 5 8 7.7975 $w=1.41688e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1735 $X2=0.2430 $Y2=0.1350
r4 5 21 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1735 $X2=0.2430 $Y2=0.2140
r5 19 20 2.85657 $w=1.3e-08 $l=1.22e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0820 $X2=0.2430 $Y2=0.0942
r6 19 18 4.37231 $w=1.3e-08 $l=1.88e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0820 $X2=0.2430 $Y2=0.0632
r7 4 8 3.2503 $w=1.53684e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1160 $X2=0.2430 $Y2=0.1350
r8 4 20 5.07188 $w=1.3e-08 $l=2.18e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1160 $X2=0.2430 $Y2=0.0942
r9 16 17 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2715
+ $Y=0.1350 $X2=0.2810 $Y2=0.1350
r10 6 16 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2615
+ $Y=0.1350 $X2=0.2715 $Y2=0.1350
r11 6 8 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2615 $Y=0.1350 $X2=0.2430 $Y2=0.1350
r12 14 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2770 $Y=0.1350
+ $X2=0.2810 $Y2=0.1350
r13 12 14 4.43042 $w=1.53e-08 $l=7.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.2845 $Y=0.1350 $X2=0.2770 $Y2=0.1350
r14 1 11 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.2885
+ $Y=0.1350 $X2=0.2985 $Y2=0.1350
r15 1 12 1.86855 $w=1.78125e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.2885 $Y=0.1350 $X2=0.2845 $Y2=0.1350
r16 3 11 2.53453 $w=1.32811e-07 $l=1.5e-09 $layer=LIG $thickness=5.23243e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2985 $Y2=0.1350
r17 3 12 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2845 $Y2=0.1350
.ends

.subckt PM_DFFHQNx2_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.00485261f
.ends

.subckt PM_DFFHQNx2_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.00416242f
.ends

.subckt PM_DFFHQNx2_ASAP7_75t_R%CLK VSS 10 3 8 5 1 6 7 4
c1 1 VSS 0.00248101f
c2 3 VSS 0.0596823f
c3 4 VSS 0.000950695f
c4 5 VSS 0.0040035f
c5 6 VSS 0.00388743f
c6 7 VSS 0.00220256f
c7 8 VSS 0.00207414f
r1 6 18 3.22357 $w=2.26279e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.2125 $X2=0.1080 $Y2=0.1820
r2 5 16 3.22357 $w=2.26279e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0575 $X2=0.1080 $Y2=0.0880
r3 17 18 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.1820 $X2=0.1080 $Y2=0.1820
r4 8 14 0.54189 $w=3.37e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1820 $X2=0.0810 $Y2=0.1630
r5 8 17 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1820 $X2=0.0945 $Y2=0.1820
r6 15 16 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.0880 $X2=0.1080 $Y2=0.0880
r7 7 15 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0880 $X2=0.0945 $Y2=0.0880
r8 13 14 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1530 $X2=0.0810 $Y2=0.1630
r9 12 13 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1530
r10 11 12 2.85657 $w=1.3e-08 $l=1.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1227 $X2=0.0810 $Y2=0.1350
r11 10 11 0.874462 $w=1.3e-08 $l=3.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1227
r12 10 4 1.57403 $w=1.3e-08 $l=6.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1122
r13 4 7 1.76614 $w=2.65738e-08 $l=2.42e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1122 $X2=0.0810 $Y2=0.0880
r14 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r15 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_DFFHQNx2_ASAP7_75t_R%PD2 VSS 7 12 4 5 1
c1 1 VSS 0.00730035f
c2 4 VSS 0.0018873f
c3 5 VSS 0.0023344f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4880 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r3 9 5 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.4605
+ $Y=0.2295 $X2=0.4860 $Y2=0.2295
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.4455
+ $Y=0.2295 $X2=0.4605 $Y2=0.2295
r5 1 8 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4320
+ $Y=0.2295 $X2=0.4455 $Y2=0.2295
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2295 $X2=0.4300 $Y2=0.2295
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2295 $X2=0.4175 $Y2=0.2295
.ends

.subckt PM_DFFHQNx2_ASAP7_75t_R%PD1 VSS 7 10 5 4 1
c1 1 VSS 0.0106263f
c2 4 VSS 0.00318954f
c3 5 VSS 0.00185362f
r1 10 9 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r2 8 9 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r3 5 8 0.123457 $w=8.1e-08 $l=1e-08 $layer=N_src_drn $thickness=1e-09 $X=0.3780
+ $Y=0.0675 $X2=0.3880 $Y2=0.0675
r4 4 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3220 $Y2=0.0675
r5 7 4 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r6 1 5 1e-05
.ends

.subckt PM_DFFHQNx2_ASAP7_75t_R%NET15 VSS 9 49 53 59 63 10 18 14 12 3 15 4 16
+ 19 17 20 1
c1 1 VSS 0.00036151f
c2 3 VSS 0.00584062f
c3 4 VSS 0.00560572f
c4 9 VSS 0.0363946f
c5 10 VSS 0.00226939f
c6 11 VSS 9.01671e-20
c7 12 VSS 0.00280457f
c8 13 VSS 6.90824e-20
c9 14 VSS 0.00883669f
c10 15 VSS 0.00138648f
c11 16 VSS 0.000721404f
c12 17 VSS 0.000428257f
c13 18 VSS 0.00607686f
c14 19 VSS 1.2124e-20
c15 20 VSS 0.00240141f
r1 63 62 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r2 61 62 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r3 3 61 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3760 $Y=0.2295 $X2=0.3880 $Y2=0.2295
r4 13 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2295 $X2=0.3760 $Y2=0.2295
r5 57 58 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r6 59 57 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.1890 $X2=0.3635 $Y2=0.1890
r7 12 58 0.185185 $w=5.4e-08 $l=1e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r8 12 3 0.518519 $w=3.9e-08 $l=4.05494e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.1890 $X2=0.3760 $Y2=0.2295
r9 3 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2295
+ $X2=0.3780 $Y2=0.2340
r10 53 52 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r11 51 52 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4420 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r12 4 51 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4300 $Y=0.0405 $X2=0.4420 $Y2=0.0405
r13 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0405 $X2=0.4300 $Y2=0.0405
r14 10 4 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0810 $X2=0.4300 $Y2=0.0810
r15 49 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0810 $X2=0.4175 $Y2=0.0810
r16 45 46 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r17 43 46 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r18 42 43 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4160
+ $Y=0.2340 $X2=0.4050 $Y2=0.2340
r19 14 20 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4340
+ $Y=0.2340 $X2=0.4590 $Y2=0.2340
r20 14 42 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4340
+ $Y=0.2340 $X2=0.4160 $Y2=0.2340
r21 4 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0405
+ $X2=0.4320 $Y2=0.0360
r22 20 34 3.01468 $w=1.741e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4590 $Y2=0.2140
r23 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4455 $Y2=0.0360
r24 18 31 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4590 $Y2=0.0630
r25 18 37 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4455 $Y2=0.0360
r26 33 34 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1850 $X2=0.4590 $Y2=0.2140
r27 32 33 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1660 $X2=0.4590 $Y2=0.1850
r28 16 19 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1525 $X2=0.4590 $Y2=0.1310
r29 16 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1525 $X2=0.4590 $Y2=0.1660
r30 30 31 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0900 $X2=0.4590 $Y2=0.0630
r31 29 30 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1025 $X2=0.4590 $Y2=0.0900
r32 15 19 2.78392 $w=1.56471e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1140 $X2=0.4590 $Y2=0.1310
r33 15 29 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1140 $X2=0.4590 $Y2=0.1025
r34 19 28 4.18306 $w=1.49565e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1310 $X2=0.4820 $Y2=0.1310
r35 27 28 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5000
+ $Y=0.1310 $X2=0.4820 $Y2=0.1310
r36 26 27 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1310 $X2=0.5000 $Y2=0.1310
r37 17 25 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1310 $X2=0.5670 $Y2=0.1310
r38 17 26 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1310 $X2=0.5130 $Y2=0.1310
r39 1 22 2.36633 $w=2.3e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.5670
+ $Y=0.1305 $X2=0.5670 $Y2=0.1305
r40 1 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1305
+ $X2=0.5670 $Y2=0.1310
r41 9 22 0.314665 $w=2.27e-07 $l=4.5e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5670 $Y=0.1350 $X2=0.5670 $Y2=0.1305
r42 3 12 1e-05
.ends

.subckt PM_DFFHQNx2_ASAP7_75t_R%noxref_26 VSS 1
c1 1 VSS 0.041505f
.ends

.subckt PM_DFFHQNx2_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.00422035f
.ends

.subckt PM_DFFHQNx2_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.00426912f
.ends

.subckt PM_DFFHQNx2_ASAP7_75t_R%NET29 VSS 10 41 44 48 50 13 17 18 14 3 15 12 1
+ 11 4 16
c1 1 VSS 0.00215637f
c2 3 VSS 0.00567591f
c3 4 VSS 0.00936239f
c4 10 VSS 0.037516f
c5 11 VSS 0.00302832f
c6 12 VSS 0.00284374f
c7 13 VSS 0.00240982f
c8 14 VSS 0.00185523f
c9 15 VSS 0.00401427f
c10 16 VSS 0.00177841f
c11 17 VSS 0.0012511f
c12 18 VSS 0.000447805f
c13 19 VSS 0.00278307f
r1 50 49 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.2295 $X2=0.6625 $Y2=0.2295
r2 13 49 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6500 $Y=0.2295 $X2=0.6625 $Y2=0.2295
r3 12 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2295 $X2=0.5920 $Y2=0.2295
r4 48 12 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.2295 $X2=0.5795 $Y2=0.2295
r5 45 13 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6210 $Y=0.2295 $X2=0.6480 $Y2=0.2295
r6 4 45 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08 $X=0.5940
+ $Y=0.2295 $X2=0.6210 $Y2=0.2295
r7 4 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2295
+ $X2=0.5940 $Y2=0.2340
r8 15 19 5.06479 $w=1.46038e-08 $l=2.70046e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5940 $Y=0.2340 $X2=0.6210 $Y2=0.2335
r9 44 43 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.0405 $X2=0.6085 $Y2=0.0405
r10 42 43 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6040 $Y=0.0405 $X2=0.6085 $Y2=0.0405
r11 3 42 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5920 $Y=0.0405 $X2=0.6040 $Y2=0.0405
r12 11 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.0405 $X2=0.5920 $Y2=0.0405
r13 41 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0405 $X2=0.5795 $Y2=0.0405
r14 19 36 0.983973 $w=1.77222e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.2335 $X2=0.6210 $Y2=0.2245
r15 3 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0405
+ $X2=0.5940 $Y2=0.0540
r16 35 36 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.2135 $X2=0.6210 $Y2=0.2245
r17 34 35 6.64591 $w=1.3e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1850 $X2=0.6210 $Y2=0.2135
r18 33 34 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1660 $X2=0.6210 $Y2=0.1850
r19 32 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1525 $X2=0.6210 $Y2=0.1660
r20 31 32 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1310 $X2=0.6210 $Y2=0.1525
r21 30 31 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1115 $X2=0.6210 $Y2=0.1310
r22 17 28 1.15159 $w=1.75e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1000 $X2=0.6210 $Y2=0.0900
r23 17 30 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1000 $X2=0.6210 $Y2=0.1115
r24 16 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0540 $X2=0.5940 $Y2=0.0720
r25 27 28 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6075 $Y=0.0900 $X2=0.6210 $Y2=0.0900
r26 18 26 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5940 $Y=0.0900 $X2=0.5805 $Y2=0.0900
r27 18 27 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5940 $Y=0.0900 $X2=0.6075 $Y2=0.0900
r28 18 29 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0900 $X2=0.5940 $Y2=0.0720
r29 25 26 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5490
+ $Y=0.0900 $X2=0.5805 $Y2=0.0900
r30 24 25 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0900 $X2=0.5490 $Y2=0.0900
r31 14 24 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5000
+ $Y=0.0900 $X2=0.5130 $Y2=0.0900
r32 1 21 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.5130
+ $Y=0.0900 $X2=0.5130 $Y2=0.0900
r33 1 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.0900
+ $X2=0.5130 $Y2=0.0900
r34 10 21 0.314665 $w=2.27e-07 $l=4.5e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5130 $Y2=0.0900
.ends

.subckt PM_DFFHQNx2_ASAP7_75t_R%PD5 VSS 7 12 4 1 5
c1 1 VSS 0.00741202f
c2 4 VSS 0.00187913f
c3 5 VSS 0.00237532f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.0405 $X2=0.7705 $Y2=0.0405
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7580 $Y=0.0405 $X2=0.7705 $Y2=0.0405
r3 9 5 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.7425
+ $Y=0.0405 $X2=0.7560 $Y2=0.0405
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.7275
+ $Y=0.0405 $X2=0.7425 $Y2=0.0405
r5 1 8 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.7020
+ $Y=0.0405 $X2=0.7275 $Y2=0.0405
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.0405 $X2=0.7000 $Y2=0.0405
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.0405 $X2=0.6875 $Y2=0.0405
.ends

.subckt PM_DFFHQNx2_ASAP7_75t_R%QN VSS 24 16 17 28 29 7 8 11 1 2
c1 1 VSS 0.00979919f
c2 2 VSS 0.0105394f
c3 7 VSS 0.00455267f
c4 8 VSS 0.00455406f
c5 9 VSS 0.0078419f
c6 10 VSS 0.00796869f
c7 11 VSS 0.00661099f
c8 12 VSS 0.00263523f
c9 13 VSS 0.00259846f
r1 29 27 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0430 $Y=0.2025 $X2=1.0405 $Y2=0.2025
r2 2 27 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0260 $Y=0.2025 $X2=1.0405 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0115 $Y=0.2025 $X2=1.0260 $Y2=0.2025
r4 28 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0090 $Y=0.2025 $X2=1.0115 $Y2=0.2025
r5 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0260 $Y=0.2025
+ $X2=1.0260 $Y2=0.2250
r6 24 25 1.69063 $w=1.3e-08 $l=7.2e-09 $layer=M1 $thickness=3.6e-08 $X=1.0850
+ $Y=0.2250 $X2=1.0922 $Y2=0.2250
r7 24 23 5.88804 $w=1.3e-08 $l=2.53e-08 $layer=M1 $thickness=3.6e-08 $X=1.0850
+ $Y=0.2250 $X2=1.0597 $Y2=0.2250
r8 22 23 7.87015 $w=1.3e-08 $l=3.37e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.2250 $X2=1.0597 $Y2=0.2250
r9 10 22 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.0145
+ $Y=0.2250 $X2=1.0260 $Y2=0.2250
r10 13 21 6.16274 $w=1.56328e-08 $l=3.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1080 $Y=0.2250 $X2=1.1080 $Y2=0.1915
r11 13 25 2.02363 $w=1.58571e-08 $l=1.58e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1080 $Y=0.2250 $X2=1.0922 $Y2=0.2250
r12 20 21 14.691 $w=1.3e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.1080
+ $Y=0.1285 $X2=1.1080 $Y2=0.1915
r13 11 12 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1080 $Y=0.0720 $X2=1.1080 $Y2=0.0450
r14 11 20 13.1752 $w=1.3e-08 $l=5.65e-08 $layer=M1 $thickness=3.6e-08 $X=1.1080
+ $Y=0.0720 $X2=1.1080 $Y2=0.1285
r15 12 19 7.91167 $w=1.40976e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1080 $Y=0.0450 $X2=1.0670 $Y2=0.0450
r16 18 19 9.56078 $w=1.3e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.0450 $X2=1.0670 $Y2=0.0450
r17 9 18 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.0145
+ $Y=0.0450 $X2=1.0260 $Y2=0.0450
r18 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0260 $Y=0.0675
+ $X2=1.0260 $Y2=0.0450
r19 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.0430 $Y=0.0675 $X2=1.0405 $Y2=0.0675
r20 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.0260 $Y=0.0675 $X2=1.0405 $Y2=0.0675
r21 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.0115 $Y=0.0675 $X2=1.0260 $Y2=0.0675
r22 16 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.0090 $Y=0.0675 $X2=1.0115 $Y2=0.0675
.ends

.subckt PM_DFFHQNx2_ASAP7_75t_R%noxref_28 VSS 1
c1 1 VSS 0.0423834f
.ends

.subckt PM_DFFHQNx2_ASAP7_75t_R%noxref_29 VSS 1
c1 1 VSS 0.0423369f
.ends

.subckt PM_DFFHQNx2_ASAP7_75t_R%noxref_27 VSS 1
c1 1 VSS 0.0415f
.ends

.subckt PM_DFFHQNx2_ASAP7_75t_R%CLKB VSS 14 15 16 17 81 83 18 20 26 6 7 23 24 4
+ 25 22 19 1 21 8 2
c1 1 VSS 0.00179184f
c2 2 VSS 0.000802772f
c3 3 VSS 0.000754022f
c4 4 VSS 0.00115302f
c5 6 VSS 0.00885416f
c6 7 VSS 0.0085707f
c7 8 VSS 0.00504283f
c8 14 VSS 0.00605314f
c9 15 VSS 0.00581477f
c10 16 VSS 0.00510025f
c11 17 VSS 0.00592939f
c12 18 VSS 0.00548094f
c13 19 VSS 0.00547471f
c14 20 VSS 0.00411307f
c15 21 VSS 0.00335428f
c16 22 VSS 0.0028383f
c17 23 VSS 0.00687114f
c18 24 VSS 0.0060817f
c19 25 VSS 0.00126875f
c20 26 VSS 0.00549311f
r1 19 7 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1600 $Y2=0.2160
r2 83 19 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r3 18 6 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1600 $Y2=0.0540
r4 81 18 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r5 4 79 2.78395 $w=2.4e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08 $X=0.7290
+ $Y=0.1780 $X2=0.7250 $Y2=0.1780
r6 17 4 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.7290 $Y=0.1350 $X2=0.7290 $Y2=0.1780
r7 3 72 10.3807 $w=2.30357e-08 $l=0 $layer=LISD $thickness=3.675e-08 $X=0.6210
+ $Y=0.1780 $X2=0.6210 $Y2=0.1780
r8 16 3 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.6210 $Y=0.1350 $X2=0.6210 $Y2=0.1780
r9 2 65 2.78395 $w=2.4e-08 $l=5e-09 $layer=LIG $thickness=4.8e-08 $X=0.4590
+ $Y=0.1780 $X2=0.4640 $Y2=0.1780
r10 15 2 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4590 $Y2=0.1780
r11 7 57 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1655 $Y2=0.2340
r12 6 53 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1655 $Y2=0.0360
r13 78 79 4.8113 $w=2.22e-08 $l=1.5e-09 $layer=LISD $thickness=2.7e-08
+ $X=0.7235 $Y=0.1780 $X2=0.7250 $Y2=0.1780
r14 77 78 10.8887 $w=2.22e-08 $l=2.15e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7020 $Y=0.1780 $X2=0.7235 $Y2=0.1780
r15 76 77 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6885 $Y=0.1780 $X2=0.7020 $Y2=0.1780
r16 75 76 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6750 $Y=0.1780 $X2=0.6885 $Y2=0.1780
r17 74 75 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6615 $Y=0.1780 $X2=0.6750 $Y2=0.1780
r18 73 74 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6480 $Y=0.1780 $X2=0.6615 $Y2=0.1780
r19 72 73 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6210 $Y=0.1780 $X2=0.6480 $Y2=0.1780
r20 71 72 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5940 $Y=0.1780 $X2=0.6210 $Y2=0.1780
r21 70 71 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5805 $Y=0.1780 $X2=0.5940 $Y2=0.1780
r22 69 70 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5670 $Y=0.1780 $X2=0.5805 $Y2=0.1780
r23 68 69 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5535 $Y=0.1780 $X2=0.5670 $Y2=0.1780
r24 67 68 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5400 $Y=0.1780 $X2=0.5535 $Y2=0.1780
r25 66 67 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5265 $Y=0.1780 $X2=0.5400 $Y2=0.1780
r26 64 65 10.3823 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4775 $Y=0.1780 $X2=0.4640 $Y2=0.1780
r27 63 64 11.142 $w=2.22e-08 $l=2.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4995 $Y=0.1780 $X2=0.4775 $Y2=0.1780
r28 62 66 1.51936 $w=2.22e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.5235
+ $Y=0.1780 $X2=0.5265 $Y2=0.1780
r29 61 62 5.31775 $w=2.22e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5130 $Y=0.1780 $X2=0.5235 $Y2=0.1780
r30 8 61 5.31775 $w=2.22e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5025 $Y=0.1780 $X2=0.5130 $Y2=0.1780
r31 8 63 1.51936 $w=2.22e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.5025
+ $Y=0.1780 $X2=0.4995 $Y2=0.1780
r32 57 58 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1655
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r33 24 50 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2340 $X2=0.1890 $Y2=0.2125
r34 24 58 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2340 $X2=0.1755 $Y2=0.2340
r35 53 54 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1655
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r36 23 49 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1890 $Y2=0.0575
r37 23 54 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1755 $Y2=0.0360
r38 51 61 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5130 $Y=0.1845
+ $X2=0.5130 $Y2=0.1780
r39 22 51 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1680 $X2=0.5130 $Y2=0.1845
r40 48 49 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0880 $X2=0.1890 $Y2=0.0575
r41 47 48 11.3097 $w=1.3e-08 $l=4.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1365 $X2=0.1890 $Y2=0.0880
r42 46 50 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1990 $X2=0.1890 $Y2=0.2125
r43 45 46 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1890 $X2=0.1890 $Y2=0.1990
r44 20 45 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1735 $X2=0.1890 $Y2=0.1890
r45 20 47 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1735 $X2=0.1890 $Y2=0.1365
r46 43 51 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.5130 $Y=0.1890
+ $X2=0.5130 $Y2=0.1845
r47 42 43 22.0364 $w=1.3e-08 $l=9.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.4185
+ $Y=0.1890 $X2=0.5130 $Y2=0.1890
r48 41 42 22.0364 $w=1.3e-08 $l=9.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1890 $X2=0.4185 $Y2=0.1890
r49 40 41 15.7403 $w=1.3e-08 $l=6.75e-08 $layer=M2 $thickness=3.6e-08 $X=0.2565
+ $Y=0.1890 $X2=0.3240 $Y2=0.1890
r50 39 40 15.7403 $w=1.3e-08 $l=6.75e-08 $layer=M2 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1890 $X2=0.2565 $Y2=0.1890
r51 39 45 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1890 $Y=0.1890
+ $X2=0.1890 $Y2=0.1890
r52 26 39 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.1775
+ $Y=0.1890 $X2=0.1890 $Y2=0.1890
r53 37 41 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.3240 $Y=0.1890
+ $X2=0.3240 $Y2=0.1890
r54 36 37 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1735 $X2=0.3240 $Y2=0.1890
r55 21 34 3.60008 $w=1.51951e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3240 $Y=0.1555 $X2=0.3240 $Y2=0.1350
r56 21 36 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1555 $X2=0.3240 $Y2=0.1735
r57 25 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r58 25 34 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3375 $Y=0.1350 $X2=0.3240 $Y2=0.1350
r59 14 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r60 1 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
.ends

.subckt PM_DFFHQNx2_ASAP7_75t_R%NET32 VSS 11 12 13 74 77 81 84 29 6 19 15 14 24
+ 17 16 18 5 26 2 23 28 27 21 22 1 25 20
c1 1 VSS 0.000782796f
c2 2 VSS 0.00812694f
c3 5 VSS 0.00501499f
c4 6 VSS 0.00494511f
c5 11 VSS 0.0374671f
c6 12 VSS 0.0809277f
c7 13 VSS 0.0809602f
c8 14 VSS 0.00504743f
c9 15 VSS 0.00526145f
c10 16 VSS 0.00910086f
c11 17 VSS 0.00197388f
c12 18 VSS 0.00185666f
c13 19 VSS 0.00276721f
c14 20 VSS 0.000821129f
c15 21 VSS 0.000535951f
c16 22 VSS 0.00142505f
c17 23 VSS 0.00383717f
c18 24 VSS 0.0062229f
c19 25 VSS 0.00233818f
c20 26 VSS 0.000131038f
c21 27 VSS 0.000406587f
c22 28 VSS 0.00038392f
c23 29 VSS 0.0113156f
r1 84 83 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r2 5 83 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6500 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r3 80 5 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6380 $Y=0.0405 $X2=0.6500 $Y2=0.0405
r4 14 80 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0405 $X2=0.6380 $Y2=0.0405
r5 81 14 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.0405 $X2=0.6335 $Y2=0.0405
r6 13 68 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=1.0530
+ $Y=0.1350 $X2=1.0530 $Y2=0.1360
r7 12 60 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.9990 $Y=0.1350 $X2=0.9990 $Y2=0.1360
r8 77 76 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r9 75 76 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7120 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r10 6 75 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7000 $Y=0.2295 $X2=0.7120 $Y2=0.2295
r11 15 6 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.2295 $X2=0.7000 $Y2=0.2295
r12 74 15 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.2295 $X2=0.6875 $Y2=0.2295
r13 5 58 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.0405
+ $X2=0.6480 $Y2=0.0360
r14 66 68 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.0405 $Y=0.1360 $X2=1.0530 $Y2=0.1360
r15 65 66 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.0260 $Y=0.1360 $X2=1.0405 $Y2=0.1360
r16 63 65 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.0115 $Y=0.1360 $X2=1.0260 $Y2=0.1360
r17 61 63 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=1.0085 $Y=0.1360 $X2=1.0115 $Y2=0.1360
r18 60 61 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.9990
+ $Y=0.1360 $X2=1.0085 $Y2=0.1360
r19 2 60 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.9895
+ $Y=0.1360 $X2=0.9990 $Y2=0.1360
r20 6 51 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7020 $Y=0.2295
+ $X2=0.7020 $Y2=0.2330
r21 58 59 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6480
+ $Y=0.0360 $X2=0.6615 $Y2=0.0360
r22 56 59 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0360 $X2=0.6615 $Y2=0.0360
r23 55 56 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6860
+ $Y=0.0360 $X2=0.6750 $Y2=0.0360
r24 16 25 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.7040
+ $Y=0.0360 $X2=0.7290 $Y2=0.0360
r25 16 55 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7040
+ $Y=0.0360 $X2=0.6860 $Y2=0.0360
r26 53 60 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.9990 $Y=0.1445
+ $X2=0.9990 $Y2=0.1360
r27 23 53 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.9990
+ $Y=0.1085 $X2=0.9990 $Y2=0.1445
r28 51 52 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.2330 $X2=0.7155 $Y2=0.2330
r29 24 52 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.2330 $X2=0.7155 $Y2=0.2330
r30 25 44 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.0360 $X2=0.7290 $Y2=0.0630
r31 48 53 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.9990 $Y=0.1530
+ $X2=0.9990 $Y2=0.1445
r32 47 48 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1530 $X2=0.9990 $Y2=0.1530
r33 46 47 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1530 $X2=0.9450 $Y2=0.1530
r34 29 46 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.8795
+ $Y=0.1530 $X2=0.8910 $Y2=0.1530
r35 45 46 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.8910 $Y=0.1485 $X2=0.8910
+ $Y2=0.1530
r36 22 45 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1305 $X2=0.8910 $Y2=0.1485
r37 18 39 6.38362 $w=1.33509e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1975 $X2=0.7290 $Y2=0.1690
r38 18 24 7.09793 $w=1.42676e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1975 $X2=0.7290 $Y2=0.2330
r39 43 44 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.0900 $X2=0.7290 $Y2=0.0630
r40 42 43 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1000 $X2=0.7290 $Y2=0.0900
r41 41 42 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1100 $X2=0.7290 $Y2=0.1000
r42 17 26 4.67854 $w=1.44583e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1360 $X2=0.7290 $Y2=0.1600
r43 17 41 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1360 $X2=0.7290 $Y2=0.1100
r44 28 40 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1575 $X2=0.8910 $Y2=0.1665
r45 28 45 1.50855 $w=1.55e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1575 $X2=0.8910 $Y2=0.1485
r46 28 46 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.8910 $Y=0.1575 $X2=0.8910
+ $Y2=0.1530
r47 26 39 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1600 $X2=0.7290 $Y2=0.1690
r48 38 40 4.19024 $w=1.156e-08 $l=2.54018e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8660 $Y=0.1620 $X2=0.8910 $Y2=0.1665
r49 21 27 1.38478 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8480 $Y=0.1620 $X2=0.8370 $Y2=0.1620
r50 21 38 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8480
+ $Y=0.1620 $X2=0.8660 $Y2=0.1620
r51 37 39 4.4015 $w=1.35e-08 $l=2.78927e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7560 $Y=0.1620 $X2=0.7290 $Y2=0.1690
r52 36 37 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1620 $X2=0.7560 $Y2=0.1620
r53 19 27 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.1620 $X2=0.8370 $Y2=0.1620
r54 19 36 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.1620 $X2=0.7830 $Y2=0.1620
r55 27 35 4.88263 $w=1.47308e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8370 $Y=0.1620 $X2=0.8370 $Y2=0.1360
r56 20 35 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1180 $X2=0.8370 $Y2=0.1360
r57 11 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.8370
+ $Y=0.1350 $X2=0.8370 $Y2=0.1350
r58 1 35 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8370 $Y=0.1350
+ $X2=0.8370 $Y2=0.1360
.ends

.subckt PM_DFFHQNx2_ASAP7_75t_R%NET37 VSS 9 32 45 12 10 11 15 4 3 14 1 16 13
c1 1 VSS 0.00103979f
c2 3 VSS 0.00624476f
c3 4 VSS 0.00663239f
c4 9 VSS 0.0384419f
c5 10 VSS 0.00329117f
c6 11 VSS 0.003282f
c7 12 VSS 0.00186966f
c8 13 VSS 0.0137838f
c9 14 VSS 0.009249f
c10 15 VSS 0.00752744f
c11 16 VSS 0.00324012f
c12 17 VSS 0.00378962f
c13 18 VSS 0.00333079f
r1 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.2295 $X2=0.8620 $Y2=0.2295
r2 45 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.2295 $X2=0.8495 $Y2=0.2295
r3 4 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.2295
+ $X2=0.8640 $Y2=0.2340
r4 42 43 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.2340 $X2=0.8865 $Y2=0.2340
r5 14 18 4.65662 $w=1.4e-08 $l=2.73724e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9180 $Y=0.2340 $X2=0.9450 $Y2=0.2295
r6 14 43 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.2340 $X2=0.8865 $Y2=0.2340
r7 18 39 0.575795 $w=1.75e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.2295 $X2=0.9450 $Y2=0.2245
r8 38 39 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.2200 $X2=0.9450 $Y2=0.2245
r9 37 38 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1935 $X2=0.9450 $Y2=0.2200
r10 36 37 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1690 $X2=0.9450 $Y2=0.1935
r11 35 36 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1420 $X2=0.9450 $Y2=0.1690
r12 34 35 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1035 $X2=0.9450 $Y2=0.1420
r13 33 34 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.0720 $X2=0.9450 $Y2=0.1035
r14 15 30 1.50855 $w=1.55e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.0495 $X2=0.9450 $Y2=0.0405
r15 15 33 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.0495 $X2=0.9450 $Y2=0.0720
r16 10 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.0405 $X2=0.8620 $Y2=0.0405
r17 32 10 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.0405 $X2=0.8495 $Y2=0.0405
r18 17 29 4.65662 $w=1.4e-08 $l=2.73724e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.0315 $X2=0.9180 $Y2=0.0360
r19 17 30 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.0315 $X2=0.9450 $Y2=0.0405
r20 3 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.0405
+ $X2=0.8640 $Y2=0.0360
r21 28 29 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.0360 $X2=0.9180 $Y2=0.0360
r22 27 28 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.0360 $X2=0.8910 $Y2=0.0360
r23 26 27 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.0360 $X2=0.8640 $Y2=0.0360
r24 13 16 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.0360 $X2=0.7830 $Y2=0.0360
r25 13 26 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0360 $X2=0.8370 $Y2=0.0360
r26 12 23 8.04505 $w=1.3e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.0705 $X2=0.7830 $Y2=0.1050
r27 12 16 6.39593 $w=1.55565e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7830 $Y=0.0705 $X2=0.7830 $Y2=0.0360
r28 1 20 2.36633 $w=2.3e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.7830
+ $Y=0.1055 $X2=0.7830 $Y2=0.1055
r29 1 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7830 $Y=0.1055
+ $X2=0.7830 $Y2=0.1050
r30 9 20 0.314665 $w=2.27e-07 $l=2.95e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.7830 $Y=0.1350 $X2=0.7830 $Y2=0.1055
.ends

.subckt PM_DFFHQNx2_ASAP7_75t_R%CLKN VSS 13 14 15 77 79 22 8 26 7 16 17 1 19 21
+ 20 18 28 23 2 24 3
c1 1 VSS 0.00161785f
c2 2 VSS 4.47588e-20
c3 3 VSS 0.000154734f
c4 7 VSS 0.0074887f
c5 8 VSS 0.00761668f
c6 13 VSS 0.0596081f
c7 14 VSS 0.00439493f
c8 15 VSS 0.0045813f
c9 16 VSS 0.00601033f
c10 17 VSS 0.00593711f
c11 18 VSS 0.00529977f
c12 19 VSS 0.00348201f
c13 20 VSS 0.00462088f
c14 21 VSS 0.00450967f
c15 22 VSS 0.000592173f
c16 23 VSS 0.000585389f
c17 24 VSS 0.00136469f
c18 25 VSS 0.0036607f
c19 26 VSS 0.00153747f
c20 27 VSS 0.00378408f
c21 28 VSS 0.0231235f
r1 79 78 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r2 17 78 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r3 77 76 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r4 16 76 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r5 8 74 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0550 $Y2=0.2340
r6 7 71 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0550 $Y2=0.0360
r7 73 74 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.2340 $X2=0.0550 $Y2=0.2340
r8 21 73 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0460 $Y2=0.2340
r9 21 27 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0180 $Y2=0.2340
r10 70 71 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.0360 $X2=0.0550 $Y2=0.0360
r11 20 70 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0460 $Y2=0.0360
r12 20 25 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0180 $Y2=0.0360
r13 27 63 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.2340 $X2=0.0180 $Y2=0.2125
r14 25 61 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.0360 $X2=0.0180 $Y2=0.0575
r15 3 58 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6750 $Y=0.1350
+ $X2=0.6750 $Y2=0.1440
r16 15 3 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6750
+ $Y=0.1350 $X2=0.6750 $Y2=0.1350
r17 2 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
r18 14 2 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r19 62 63 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1820 $X2=0.0180 $Y2=0.2125
r20 19 26 0.998523 $w=1.74118e-08 $l=1.01119e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1630 $X2=0.0165 $Y2=0.1530
r21 19 62 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1630 $X2=0.0180 $Y2=0.1820
r22 60 61 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0880 $X2=0.0180 $Y2=0.0575
r23 18 26 5.19594 $w=1.44151e-08 $l=2.80401e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1250 $X2=0.0165 $Y2=0.1530
r24 18 60 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1250 $X2=0.0180 $Y2=0.0880
r25 24 58 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1135 $X2=0.6750 $Y2=0.1440
r26 23 56 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1530
r27 52 53 1.90199 $w=1.38333e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.0255 $Y=0.1530 $X2=0.0345 $Y2=0.1530
r28 26 52 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0165
+ $Y=0.1530 $X2=0.0255 $Y2=0.1530
r29 50 58 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.6750 $Y=0.1530
+ $X2=0.6750 $Y2=0.1440
r30 49 50 18.3054 $w=1.3e-08 $l=7.85e-08 $layer=M2 $thickness=3.6e-08 $X=0.5965
+ $Y=0.1530 $X2=0.6750 $Y2=0.1530
r31 48 49 29.3819 $w=1.3e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.4705
+ $Y=0.1530 $X2=0.5965 $Y2=0.1530
r32 47 48 15.2739 $w=1.3e-08 $l=6.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1530 $X2=0.4705 $Y2=0.1530
r33 47 56 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4050 $Y=0.1530
+ $X2=0.4050 $Y2=0.1530
r34 46 47 27.8662 $w=1.3e-08 $l=1.195e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.2855 $Y=0.1530 $X2=0.4050 $Y2=0.1530
r35 45 46 27.5164 $w=1.3e-08 $l=1.18e-07 $layer=M2 $thickness=3.6e-08 $X=0.1675
+ $Y=0.1530 $X2=0.2855 $Y2=0.1530
r36 44 45 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M2 $thickness=3.6e-08 $X=0.1510
+ $Y=0.1530 $X2=0.1675 $Y2=0.1530
r37 43 44 13.7582 $w=1.3e-08 $l=5.9e-08 $layer=M2 $thickness=3.6e-08 $X=0.0920
+ $Y=0.1530 $X2=0.1510 $Y2=0.1530
r38 42 43 13.7582 $w=1.3e-08 $l=5.9e-08 $layer=M2 $thickness=3.6e-08 $X=0.0330
+ $Y=0.1530 $X2=0.0920 $Y2=0.1530
r39 42 53 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.0330 $Y=0.1530
+ $X2=0.0345 $Y2=0.1530
r40 28 42 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.0215
+ $Y=0.1530 $X2=0.0330 $Y2=0.1530
r41 39 44 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1510 $Y=0.1440
+ $X2=0.1510 $Y2=0.1530
r42 22 39 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1510
+ $Y=0.1160 $X2=0.1510 $Y2=0.1440
r43 37 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1550 $Y=0.1350
+ $X2=0.1510 $Y2=0.1440
r44 36 37 4.43042 $w=1.53e-08 $l=7.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1475 $Y=0.1350 $X2=0.1550 $Y2=0.1350
r45 34 36 1.86855 $w=1.78125e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1435 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r46 1 34 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.1335
+ $Y=0.1350 $X2=0.1435 $Y2=0.1350
r47 13 1 2.53453 $w=1.32811e-07 $l=1.5e-09 $layer=LIG $thickness=5.23243e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1335 $Y2=0.1350
r48 13 36 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r49 8 17 1e-05
r50 7 16 1e-05
.ends


*
.SUBCKT DFFHQNx2_ASAP7_75t_R VSS VDD CLK D QN
*
* VSS VSS
* VDD VDD
* CLK CLK
* D D
* QN QN
*
*

MM20 N_MM20_d N_MM20_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM23 N_MM23_d N_MM22_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM10_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM6 N_MM6_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM12 N_MM12_d N_MM12_g N_MM12_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM17 N_MM17_d N_MM13_g N_MM17_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM16 N_MM16_d N_MM19_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM14 N_MM14_d N_MM14_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM24 N_MM24_d N_MM24_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@2 N_MM24@2_d N_MM24@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM21 N_MM21_d N_MM20_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM22 N_MM22_d N_MM22_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM13 N_MM13_d N_MM13_g N_MM13_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM18 N_MM18_d N_MM18_g N_MM18_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM19 N_MM19_d N_MM19_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM15 N_MM15_d N_MM14_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM25 N_MM25_d N_MM24_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@2 N_MM25@2_d N_MM24@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "DFFHQNx2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "DFFHQNx2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_DFFHQNx2_ASAP7_75t_R%PD3 VSS N_MM9_s N_MM8_d N_PD3_1
+ PM_DFFHQNx2_ASAP7_75t_R%PD3
cc_1 N_PD3_1 N_MM9_g 0.00773019f
cc_2 N_PD3_1 N_MM11_g 0.00773412f
x_PM_DFFHQNx2_ASAP7_75t_R%PU1 VSS N_MM3_d N_MM1_s N_PU1_1
+ PM_DFFHQNx2_ASAP7_75t_R%PU1
cc_3 N_PU1_1 N_MM3_g 0.0171044f
cc_4 N_PU1_1 N_MM1_g 0.0169736f
x_PM_DFFHQNx2_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_DFFHQNx2_ASAP7_75t_R%noxref_23
cc_5 N_noxref_23_1 N_MM3_g 0.0018531f
cc_6 N_noxref_23_1 N_CLKB_7 0.000100589f
cc_7 N_noxref_23_1 N_CLKB_19 0.000556653f
cc_8 N_noxref_23_1 N_noxref_20_1 0.000463245f
cc_9 N_noxref_23_1 N_noxref_21_1 0.00768971f
cc_10 N_noxref_23_1 N_noxref_22_1 0.00122255f
x_PM_DFFHQNx2_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_DFFHQNx2_ASAP7_75t_R%noxref_22
cc_11 N_noxref_22_1 N_MM3_g 0.00183891f
cc_12 N_noxref_22_1 N_CLKB_6 0.000104326f
cc_13 N_noxref_22_1 N_CLKB_18 0.00055486f
cc_14 N_noxref_22_1 N_noxref_20_1 0.00768744f
cc_15 N_noxref_22_1 N_noxref_21_1 0.000463741f
x_PM_DFFHQNx2_ASAP7_75t_R%PD4 VSS N_MM18_s N_MM19_d N_PD4_1
+ PM_DFFHQNx2_ASAP7_75t_R%PD4
cc_16 N_PD4_1 N_MM18_g 0.00773071f
cc_17 N_PD4_1 N_MM19_g 0.00776505f
x_PM_DFFHQNx2_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_DFFHQNx2_ASAP7_75t_R%noxref_18
cc_18 N_noxref_18_1 N_MM20_g 0.00368318f
cc_19 N_noxref_18_1 N_CLKN_19 6.24201e-20
cc_20 N_noxref_18_1 N_CLKN_18 0.000312904f
cc_21 N_noxref_18_1 N_CLKN_7 0.000503374f
cc_22 N_noxref_18_1 N_CLKN_16 0.0278236f
x_PM_DFFHQNx2_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_DFFHQNx2_ASAP7_75t_R%noxref_21
cc_23 N_noxref_21_1 N_CLKN_1 0.000396541f
cc_24 N_noxref_21_1 N_MM22_g 0.00344681f
cc_25 N_noxref_21_1 N_CLKB_7 0.000426471f
cc_26 N_noxref_21_1 N_CLKB_19 0.0270308f
cc_27 N_noxref_21_1 N_noxref_20_1 0.00141787f
x_PM_DFFHQNx2_ASAP7_75t_R%D VSS D N_MM3_g N_D_5 N_D_6 N_D_7 N_D_9 N_D_1 N_D_4
+ N_D_8 PM_DFFHQNx2_ASAP7_75t_R%D
cc_28 N_D_5 N_CLKN_22 0.000146036f
cc_29 N_D_5 N_CLKN_23 7.47542e-20
cc_30 N_D_5 N_CLKN_1 0.000102901f
cc_31 N_D_6 N_CLKN_28 0.000654702f
cc_32 N_D_5 N_CLKN_28 0.00330841f
x_PM_DFFHQNx2_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_DFFHQNx2_ASAP7_75t_R%noxref_20
cc_33 N_noxref_20_1 N_CLKN_1 0.000398066f
cc_34 N_noxref_20_1 N_MM22_g 0.00343386f
cc_35 N_noxref_20_1 N_CLKB_6 0.000423111f
cc_36 N_noxref_20_1 N_CLKB_18 0.0270309f
x_PM_DFFHQNx2_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_DFFHQNx2_ASAP7_75t_R%noxref_19
cc_37 N_noxref_19_1 N_MM20_g 0.00367249f
cc_38 N_noxref_19_1 N_CLKN_26 8.87656e-20
cc_39 N_noxref_19_1 N_CLKN_18 0.000152591f
cc_40 N_noxref_19_1 N_CLKN_19 0.000196778f
cc_41 N_noxref_19_1 N_CLKN_8 0.000505002f
cc_42 N_noxref_19_1 N_CLKN_17 0.027853f
cc_43 N_noxref_19_1 N_noxref_18_1 0.00204786f
x_PM_DFFHQNx2_ASAP7_75t_R%CLK VSS CLK N_MM20_g N_CLK_8 N_CLK_5 N_CLK_1 N_CLK_6
+ N_CLK_7 N_CLK_4 PM_DFFHQNx2_ASAP7_75t_R%CLK
x_PM_DFFHQNx2_ASAP7_75t_R%PD2 VSS N_MM10_s N_MM11_d N_PD2_4 N_PD2_5 N_PD2_1
+ PM_DFFHQNx2_ASAP7_75t_R%PD2
cc_44 N_PD2_4 N_MM10_g 0.0150485f
cc_45 N_PD2_5 N_CLKB_8 0.00146961f
cc_46 N_PD2_1 N_CLKB_2 0.000539912f
cc_47 N_PD2_1 N_MM9_g 0.00206219f
cc_48 N_PD2_4 N_MM9_g 0.00714092f
cc_49 N_PD2_5 N_MM9_g 0.0240569f
cc_50 N_PD2_5 N_MM11_g 0.0146029f
cc_51 N_PD2_1 N_NET15_14 0.000435678f
cc_52 N_PD2_4 N_NET15_3 0.000614551f
cc_53 N_PD2_1 N_NET15_20 0.00320687f
x_PM_DFFHQNx2_ASAP7_75t_R%PD1 VSS N_MM5_d N_MM4_s N_PD1_5 N_PD1_4 N_PD1_1
+ PM_DFFHQNx2_ASAP7_75t_R%PD1
cc_54 N_PD1_5 N_CLKN_2 0.000858363f
cc_55 N_PD1_5 N_CLKN_23 0.000316649f
cc_56 N_PD1_5 N_MM10_g 0.0343214f
cc_57 N_PD1_4 N_MM3_g 0.0359359f
cc_58 N_PD1_5 N_CLKB_25 0.000413006f
cc_59 N_PD1_5 N_CLKB_1 0.00234469f
cc_60 N_PD1_5 N_MM1_g 0.0735635f
cc_61 N_PD1_1 N_NET15_4 0.0012224f
cc_62 N_PD1_1 N_NET15_10 0.00350016f
x_PM_DFFHQNx2_ASAP7_75t_R%NET15 VSS N_MM7_g N_MM4_d N_MM9_d N_MM1_d N_MM10_d
+ N_NET15_10 N_NET15_18 N_NET15_14 N_NET15_12 N_NET15_3 N_NET15_15 N_NET15_4
+ N_NET15_16 N_NET15_19 N_NET15_17 N_NET15_20 N_NET15_1
+ PM_DFFHQNx2_ASAP7_75t_R%NET15
cc_63 N_NET15_10 N_CLKN_3 0.000103938f
cc_64 N_NET15_10 N_CLKN_28 0.000104536f
cc_65 N_NET15_10 N_MM13_g 0.000188967f
cc_66 N_NET15_10 N_CLKN_23 0.000326582f
cc_67 N_NET15_18 N_CLKN_23 0.000369739f
cc_68 N_NET15_14 N_CLKN_23 0.000396037f
cc_69 N_NET15_12 N_MM10_g 0.0164257f
cc_70 N_NET15_3 N_CLKN_2 0.000773789f
cc_71 N_NET15_15 N_CLKN_23 0.00110463f
cc_72 N_NET15_4 N_MM10_g 0.00111964f
cc_73 N_NET15_3 N_MM10_g 0.0012324f
cc_74 N_NET15_16 N_CLKN_23 0.00124348f
cc_75 N_NET15_10 N_CLKN_2 0.0016475f
cc_76 N_NET15_19 N_CLKN_23 0.00296637f
cc_77 N_NET15_17 N_CLKN_28 0.00351688f
cc_78 N_NET15_10 N_MM10_g 0.0529705f
cc_79 N_NET15_10 N_CLKB_22 0.000366011f
cc_80 N_NET15_10 N_MM1_g 0.000402233f
cc_81 N_NET15_10 N_CLKB_21 0.000176977f
cc_82 N_NET15_10 N_CLKB_25 0.000272629f
cc_83 N_NET15_20 N_CLKB_22 0.000316176f
cc_84 N_NET15_16 N_CLKB_22 0.00266707f
cc_85 N_NET15_3 N_CLKB_1 0.000338008f
cc_86 N_NET15_17 N_CLKB_8 0.000557344f
cc_87 N_NET15_4 N_MM9_g 0.000623527f
cc_88 N_NET15_3 N_CLKB_21 0.000652452f
cc_89 N_NET15_1 N_CLKB_8 0.00227386f
cc_90 N_NET15_16 N_CLKB_2 0.000779279f
cc_91 N_NET15_12 N_CLKB_1 0.000794611f
cc_92 N_NET15_3 N_MM1_g 0.00175458f
cc_93 N_NET15_14 N_CLKB_26 0.00280164f
cc_94 N_NET15_17 N_CLKB_22 0.00357979f
cc_95 N_MM7_g N_CLKB_8 0.00464846f
cc_96 N_NET15_12 N_MM1_g 0.0336984f
cc_97 N_MM7_g N_MM12_g 0.0127429f
cc_98 N_NET15_10 N_MM9_g 0.0364088f
cc_99 N_NET15_17 N_MM11_g 0.000358889f
cc_100 N_NET15_4 N_NET29_1 0.000395733f
cc_101 N_NET15_17 N_NET29_1 0.000829739f
cc_102 N_MM7_g N_NET29_3 0.000906652f
cc_103 N_NET15_1 N_NET29_14 0.000924813f
cc_104 N_NET15_17 N_NET29_17 0.00101631f
cc_105 N_NET15_1 N_MM11_g 0.00114171f
cc_106 N_MM7_g N_NET29_1 0.00116102f
cc_107 N_NET15_15 N_NET29_14 0.00124193f
cc_108 N_MM7_g N_NET29_12 0.00639303f
cc_109 N_MM7_g N_NET29_11 0.00641111f
cc_110 N_NET15_17 N_NET29_14 0.00738558f
cc_111 N_MM7_g N_MM11_g 0.029375f
x_PM_DFFHQNx2_ASAP7_75t_R%noxref_26 VSS N_noxref_26_1
+ PM_DFFHQNx2_ASAP7_75t_R%noxref_26
cc_112 N_noxref_26_1 N_NET37_10 0.000646603f
cc_113 N_noxref_26_1 N_MM24_g 0.00169808f
cc_114 N_noxref_26_1 N_noxref_24_1 0.00776813f
cc_115 N_noxref_26_1 N_noxref_25_1 0.000476405f
x_PM_DFFHQNx2_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_DFFHQNx2_ASAP7_75t_R%noxref_24
cc_116 N_noxref_24_1 N_NET37_10 0.0170334f
cc_117 N_noxref_24_1 N_NET32_1 0.000196229f
cc_118 N_noxref_24_1 N_MM14_g 0.00594013f
x_PM_DFFHQNx2_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_DFFHQNx2_ASAP7_75t_R%noxref_25
cc_119 N_noxref_25_1 N_NET37_11 0.0169143f
cc_120 N_noxref_25_1 N_NET32_1 0.000200836f
cc_121 N_noxref_25_1 N_MM14_g 0.00603245f
cc_122 N_noxref_25_1 N_noxref_24_1 0.0015414f
x_PM_DFFHQNx2_ASAP7_75t_R%NET29 VSS N_MM11_g N_MM6_d N_MM12_d N_MM7_d N_MM13_d
+ N_NET29_13 N_NET29_17 N_NET29_18 N_NET29_14 N_NET29_3 N_NET29_15 N_NET29_12
+ N_NET29_1 N_NET29_11 N_NET29_4 N_NET29_16 PM_DFFHQNx2_ASAP7_75t_R%NET29
cc_123 N_NET29_13 N_MM10_g 0.000130138f
cc_124 N_NET29_13 N_CLKN_24 0.000324225f
cc_125 N_NET29_13 N_CLKN_28 0.00022929f
cc_126 N_NET29_13 N_CLKN_3 0.000229581f
cc_127 N_NET29_17 N_CLKN_24 0.00452728f
cc_128 N_NET29_17 N_CLKN_3 0.000282384f
cc_129 N_NET29_18 N_CLKN_24 0.000632715f
cc_130 N_NET29_14 N_CLKN_28 0.00279064f
cc_131 N_NET29_13 N_MM13_g 0.0153408f
cc_132 N_NET29_3 N_CLKB_8 0.00055579f
cc_133 N_NET29_3 N_CLKB_2 0.000123737f
cc_134 N_NET29_3 N_CLKB_22 0.000157982f
cc_135 N_NET29_3 N_MM9_g 0.000165533f
cc_136 N_NET29_3 N_CLKB_26 0.000172194f
cc_137 N_NET29_15 N_CLKB_22 0.000290783f
cc_138 N_NET29_12 N_MM12_g 0.0078041f
cc_139 N_NET29_13 N_MM12_g 0.00777346f
cc_140 N_NET29_15 N_CLKB_8 0.000383383f
cc_141 N_NET29_1 N_MM9_g 0.000560232f
cc_142 N_NET29_17 N_CLKB_8 0.00157509f
cc_143 N_NET29_11 N_MM12_g 0.00651789f
cc_144 N_NET29_4 N_MM12_g 0.00255242f
cc_145 N_NET29_4 N_CLKB_8 0.00635858f
cc_146 N_MM11_g N_MM9_g 0.0142053f
cc_147 N_NET29_3 N_MM12_g 0.0259349f
x_PM_DFFHQNx2_ASAP7_75t_R%PD5 VSS N_MM17_s N_MM16_d N_PD5_4 N_PD5_1 N_PD5_5
+ PM_DFFHQNx2_ASAP7_75t_R%PD5
cc_148 N_PD5_4 N_MM13_g 0.0152681f
cc_149 N_PD5_1 N_MM18_g 0.000759305f
cc_150 N_PD5_4 N_MM18_g 0.0069504f
cc_151 N_PD5_5 N_MM18_g 0.0239792f
cc_152 N_PD5_1 N_MM19_g 0.000915839f
cc_153 N_PD5_5 N_MM19_g 0.0155378f
cc_154 N_PD5_1 N_NET32_14 0.000516191f
cc_155 N_PD5_1 N_NET32_16 0.000436854f
cc_156 N_PD5_1 N_NET32_17 0.000599516f
cc_157 N_PD5_4 N_NET32_5 0.000664268f
cc_158 N_PD5_1 N_NET32_25 0.00239266f
x_PM_DFFHQNx2_ASAP7_75t_R%QN VSS QN N_MM24_d N_MM24@2_d N_MM25_d N_MM25@2_d
+ N_QN_7 N_QN_8 N_QN_11 N_QN_1 N_QN_2 PM_DFFHQNx2_ASAP7_75t_R%QN
cc_159 N_QN_7 N_NET32_23 0.00191833f
cc_160 N_QN_7 N_NET32_2 0.000491627f
cc_161 N_QN_7 N_NET32_29 0.000747871f
cc_162 N_QN_8 N_MM24@2_g 0.0309015f
cc_163 N_QN_11 N_NET32_2 0.00111203f
cc_164 N_QN_1 N_NET32_23 0.00184027f
cc_165 N_QN_1 N_MM24@2_g 0.00200269f
cc_166 N_QN_2 N_MM24@2_g 0.00214521f
cc_167 N_QN_8 N_NET32_2 0.0046795f
cc_168 N_QN_7 N_MM24_g 0.0371494f
cc_169 N_QN_7 N_MM24@2_g 0.0683592f
x_PM_DFFHQNx2_ASAP7_75t_R%noxref_28 VSS N_noxref_28_1
+ PM_DFFHQNx2_ASAP7_75t_R%noxref_28
cc_170 N_noxref_28_1 N_MM24@2_g 0.0014729f
cc_171 N_noxref_28_1 N_QN_7 0.00082904f
x_PM_DFFHQNx2_ASAP7_75t_R%noxref_29 VSS N_noxref_29_1
+ PM_DFFHQNx2_ASAP7_75t_R%noxref_29
cc_172 N_noxref_29_1 N_MM24@2_g 0.00147248f
cc_173 N_noxref_29_1 N_QN_8 0.000830971f
cc_174 N_noxref_29_1 N_noxref_28_1 0.00176864f
x_PM_DFFHQNx2_ASAP7_75t_R%noxref_27 VSS N_noxref_27_1
+ PM_DFFHQNx2_ASAP7_75t_R%noxref_27
cc_175 N_noxref_27_1 N_NET37_11 0.000632999f
cc_176 N_noxref_27_1 N_MM24_g 0.00171331f
cc_177 N_noxref_27_1 N_noxref_24_1 0.000478341f
cc_178 N_noxref_27_1 N_noxref_25_1 0.0077709f
cc_179 N_noxref_27_1 N_noxref_26_1 0.00123966f
x_PM_DFFHQNx2_ASAP7_75t_R%CLKB VSS N_MM1_g N_MM9_g N_MM12_g N_MM18_g N_MM23_d
+ N_MM22_d N_CLKB_18 N_CLKB_20 N_CLKB_26 N_CLKB_6 N_CLKB_7 N_CLKB_23 N_CLKB_24
+ N_CLKB_4 N_CLKB_25 N_CLKB_22 N_CLKB_19 N_CLKB_1 N_CLKB_21 N_CLKB_8 N_CLKB_2
+ PM_DFFHQNx2_ASAP7_75t_R%CLKB
cc_180 N_CLKB_18 N_CLK_6 8.57854e-20
cc_181 N_CLKB_20 N_CLK_6 9.12674e-20
cc_182 N_CLKB_26 N_CLK_6 0.000123346f
cc_183 N_CLKB_6 N_CLK_6 0.000361693f
cc_184 N_CLKB_7 N_CLK_6 0.000387298f
cc_185 N_CLKB_23 N_CLK_7 0.000500038f
cc_186 N_CLKB_20 N_CLK_8 0.000514673f
cc_187 N_CLKB_23 N_CLK_5 0.00120151f
cc_188 N_CLKB_24 N_CLK_6 0.00199622f
cc_189 N_CLKB_6 N_MM22_g 0.000721222f
cc_190 N_CLKB_7 N_MM22_g 0.000747071f
cc_191 N_CLKB_4 N_MM13_g 0.000222558f
cc_192 N_CLKB_25 N_CLKN_28 0.000285919f
cc_193 N_CLKB_22 N_CLKN_28 0.000669652f
cc_194 N_CLKB_24 N_CLKN_22 0.000310766f
cc_195 N_CLKB_19 N_MM22_g 0.0110945f
cc_196 N_CLKB_23 N_CLKN_22 0.000357496f
cc_197 N_CLKB_1 N_CLKN_2 0.00169517f
cc_198 N_CLKB_21 N_CLKN_28 0.00104596f
cc_199 N_CLKB_20 N_CLKN_22 0.00766617f
cc_200 N_CLKB_20 N_CLKN_28 0.000519084f
cc_201 N_CLKB_8 N_CLKN_24 0.000534456f
cc_202 N_CLKB_25 N_CLKN_2 0.000549016f
cc_203 N_CLKB_2 N_MM10_g 0.000589093f
cc_204 N_CLKB_26 N_CLKN_23 0.000616959f
cc_205 N_CLKB_8 N_CLKN_3 0.00279616f
cc_206 N_CLKB_20 N_CLKN_1 0.000691464f
cc_207 N_CLKB_19 N_CLKN_1 0.00121517f
cc_208 N_MM1_g N_MM10_g 0.0016376f
cc_209 N_CLKB_25 N_CLKN_23 0.00263609f
cc_210 N_CLKB_8 N_MM13_g 0.00423843f
cc_211 N_MM12_g N_MM13_g 0.0057228f
cc_212 N_MM9_g N_MM10_g 0.00910614f
cc_213 N_MM18_g N_MM13_g 0.0184455f
cc_214 N_CLKB_26 N_CLKN_28 0.0306393f
cc_215 N_CLKB_18 N_MM22_g 0.0388995f
cc_216 N_CLKB_6 N_MM3_g 0.00011685f
cc_217 N_CLKB_21 N_MM3_g 0.000132909f
cc_218 N_CLKB_20 N_MM3_g 0.000186961f
cc_219 N_CLKB_1 N_MM3_g 0.000265584f
cc_220 N_CLKB_25 N_MM3_g 0.000617636f
cc_221 N_CLKB_23 N_D_7 0.000854422f
cc_222 N_CLKB_26 N_D_6 0.00108917f
cc_223 N_CLKB_21 N_D_6 0.0011142f
cc_224 N_CLKB_24 N_D_9 0.00121817f
cc_225 N_CLKB_1 N_D_1 0.00161854f
cc_226 N_CLKB_20 N_D_4 0.00181181f
cc_227 N_CLKB_25 N_D_6 0.00203563f
cc_228 N_CLKB_20 N_D_5 0.00266241f
cc_229 N_CLKB_20 N_D_8 0.00411739f
cc_230 N_MM1_g N_MM3_g 0.0052732f
x_PM_DFFHQNx2_ASAP7_75t_R%NET32 VSS N_MM14_g N_MM24_g N_MM24@2_g N_MM13_s
+ N_MM18_d N_MM12_s N_MM17_d N_NET32_29 N_NET32_6 N_NET32_19 N_NET32_15
+ N_NET32_14 N_NET32_24 N_NET32_17 N_NET32_16 N_NET32_18 N_NET32_5 N_NET32_26
+ N_NET32_2 N_NET32_23 N_NET32_28 N_NET32_27 N_NET32_21 N_NET32_22 N_NET32_1
+ N_NET32_25 N_NET32_20 PM_DFFHQNx2_ASAP7_75t_R%NET32
cc_231 N_NET32_29 N_CLKN_28 0.000145615f
cc_232 N_NET32_6 N_MM13_g 0.000163831f
cc_233 N_NET32_19 N_CLKN_24 0.000218115f
cc_234 N_NET32_15 N_MM13_g 0.00675259f
cc_235 N_NET32_14 N_MM13_g 0.0067885f
cc_236 N_NET32_24 N_CLKN_24 0.000353816f
cc_237 N_NET32_17 N_CLKN_24 0.00434135f
cc_238 N_NET32_17 N_CLKN_3 0.000445115f
cc_239 N_NET32_16 N_CLKN_24 0.000508134f
cc_240 N_NET32_18 N_CLKN_24 0.000522964f
cc_241 N_NET32_5 N_CLKN_3 0.000536728f
cc_242 N_NET32_26 N_CLKN_24 0.000548919f
cc_243 N_NET32_16 N_CLKN_28 0.00107634f
cc_244 N_NET32_5 N_MM13_g 0.018421f
cc_245 N_NET32_15 N_CLKB_26 8.96432e-20
cc_246 N_NET32_24 N_CLKB_8 0.000184612f
cc_247 N_NET32_26 N_CLKB_8 0.000201135f
cc_248 N_NET32_14 N_MM12_g 0.00677653f
cc_249 N_NET32_6 N_CLKB_8 0.000297547f
cc_250 N_NET32_19 N_CLKB_4 0.000390105f
cc_251 N_NET32_17 N_CLKB_8 0.000424013f
cc_252 N_NET32_18 N_CLKB_8 0.000613378f
cc_253 N_NET32_15 N_CLKB_4 0.000928311f
cc_254 N_NET32_6 N_MM18_g 0.000989101f
cc_255 N_NET32_15 N_CLKB_8 0.00230339f
cc_256 N_NET32_5 N_MM12_g 0.00951489f
cc_257 N_NET32_15 N_MM18_g 0.0162711f
cc_258 N_NET32_17 N_NET29_3 0.000120104f
cc_259 N_NET32_24 N_NET29_3 0.00013281f
cc_260 N_NET32_6 N_NET29_3 0.000211236f
cc_261 N_NET32_15 N_NET29_3 0.000438565f
cc_262 N_NET32_14 N_NET29_3 0.000463915f
cc_263 N_NET32_24 N_NET29_4 0.000318287f
cc_264 N_NET32_6 N_NET29_4 0.000418085f
cc_265 N_NET32_16 N_NET29_16 0.000525166f
cc_266 N_NET32_15 N_NET29_4 0.000582695f
cc_267 N_NET32_24 N_NET29_17 0.000615677f
cc_268 N_NET32_16 N_NET29_18 0.00164128f
cc_269 N_NET32_5 N_NET29_3 0.00379032f
cc_270 N_NET32_16 N_MM19_g 9.65726e-20
cc_271 N_NET32_18 N_MM19_g 0.000139988f
cc_272 N_NET32_2 N_MM19_g 0.000149985f
cc_273 N_NET32_23 N_MM19_g 0.000158903f
cc_274 N_NET32_28 N_MM19_g 0.00019082f
cc_275 N_NET32_27 N_NET37_12 0.000215496f
cc_276 N_MM14_g N_NET37_10 0.00686462f
cc_277 N_MM14_g N_NET37_11 0.00682944f
cc_278 N_NET32_2 N_NET37_15 0.000267362f
cc_279 N_NET32_23 N_NET37_15 0.007259f
cc_280 N_NET32_21 N_NET37_4 0.000330589f
cc_281 N_MM14_g N_NET37_3 0.000397637f
cc_282 N_NET32_22 N_NET37_15 0.00186261f
cc_283 N_MM14_g N_NET37_4 0.000516529f
cc_284 N_NET32_21 N_NET37_14 0.000650478f
cc_285 N_NET32_1 N_NET37_1 0.000686419f
cc_286 N_NET32_25 N_NET37_16 0.000794357f
cc_287 N_NET32_17 N_NET37_1 0.000849146f
cc_288 N_NET32_28 N_NET37_15 0.00090017f
cc_289 N_NET32_20 N_NET37_12 0.000940696f
cc_290 N_NET32_22 N_NET37_13 0.00110495f
cc_291 N_MM14_g N_NET37_1 0.00113556f
cc_292 N_NET32_28 N_NET37_14 0.00127828f
cc_293 N_NET32_1 N_MM19_g 0.00129556f
cc_294 N_NET32_19 N_NET37_12 0.00153111f
cc_295 N_NET32_29 N_NET37_15 0.00187315f
cc_296 N_NET32_17 N_NET37_12 0.00471844f
cc_297 N_MM14_g N_MM19_g 0.0293451f
x_PM_DFFHQNx2_ASAP7_75t_R%NET37 VSS N_MM19_g N_MM14_d N_MM15_d N_NET37_12
+ N_NET37_10 N_NET37_11 N_NET37_15 N_NET37_4 N_NET37_3 N_NET37_14 N_NET37_1
+ N_NET37_16 N_NET37_13 PM_DFFHQNx2_ASAP7_75t_R%NET37
cc_298 N_MM19_g N_CLKB_8 0.000215376f
cc_299 N_MM19_g N_CLKB_4 0.000537906f
cc_300 N_MM19_g N_MM18_g 0.0135387f
x_PM_DFFHQNx2_ASAP7_75t_R%CLKN VSS N_MM22_g N_MM10_g N_MM13_g N_MM20_d N_MM21_d
+ N_CLKN_22 N_CLKN_8 N_CLKN_26 N_CLKN_7 N_CLKN_16 N_CLKN_17 N_CLKN_1 N_CLKN_19
+ N_CLKN_21 N_CLKN_20 N_CLKN_18 N_CLKN_28 N_CLKN_23 N_CLKN_2 N_CLKN_24 N_CLKN_3
+ PM_DFFHQNx2_ASAP7_75t_R%CLKN
cc_301 N_CLKN_22 N_MM20_g 0.000243475f
cc_302 N_CLKN_8 N_MM20_g 0.00112888f
cc_303 N_CLKN_26 N_MM20_g 0.000251231f
cc_304 N_CLKN_7 N_MM20_g 0.0011647f
cc_305 N_CLKN_16 N_MM20_g 0.0112193f
cc_306 N_CLKN_17 N_MM20_g 0.0113277f
cc_307 N_CLKN_1 N_CLK_8 0.000441582f
cc_308 N_CLKN_19 N_CLK_8 0.000504441f
cc_309 N_CLKN_21 N_CLK_8 0.000765329f
cc_310 N_CLKN_20 N_CLK_5 0.000800078f
cc_311 N_CLKN_26 N_CLK_1 0.000803931f
cc_312 N_CLKN_21 N_CLK_6 0.000842599f
cc_313 N_CLKN_22 N_CLK_7 0.001063f
cc_314 N_CLKN_18 N_CLK_7 0.00116296f
cc_315 N_CLKN_28 N_CLK_8 0.00176828f
cc_316 N_CLKN_26 N_CLK_8 0.00178252f
cc_317 N_CLKN_1 N_CLK_1 0.00248534f
cc_318 N_CLKN_20 N_CLK_7 0.00268142f
cc_319 N_CLKN_22 N_CLK_8 0.00324624f
cc_320 N_CLKN_26 N_CLK_4 0.00343261f
cc_321 N_MM22_g N_MM20_g 0.0350536f
*END of DFFHQNx2_ASAP7_75t_R.pxi
.ENDS
** Design:	DFFHQNx3_ASAP7_75t_R
* Created:	"Fri Aug 17 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "DFFHQNx3_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "DFFHQNx3_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_DFFHQNx3_ASAP7_75t_R%noxref_27 VSS 1
c1 1 VSS 0.0414884f
.ends

.subckt PM_DFFHQNx3_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.00423187f
.ends

.subckt PM_DFFHQNx3_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.00427325f
.ends

.subckt PM_DFFHQNx3_ASAP7_75t_R%noxref_29 VSS 1
c1 1 VSS 0.00530902f
.ends

.subckt PM_DFFHQNx3_ASAP7_75t_R%noxref_28 VSS 1
c1 1 VSS 0.00558735f
.ends

.subckt PM_DFFHQNx3_ASAP7_75t_R%noxref_26 VSS 1
c1 1 VSS 0.0414956f
.ends

.subckt PM_DFFHQNx3_ASAP7_75t_R%QN VSS 31 24 25 35 42 43 45 13 19 18 15 3 4 2 1
+ 16 14
c1 1 VSS 0.0104295f
c2 2 VSS 0.0114933f
c3 3 VSS 0.00800468f
c4 4 VSS 0.00789496f
c5 13 VSS 0.00455675f
c6 14 VSS 0.00343097f
c7 15 VSS 0.00455816f
c8 16 VSS 0.00344889f
c9 17 VSS 0.0148664f
c10 18 VSS 0.014522f
c11 19 VSS 0.00377841f
c12 20 VSS 0.00271351f
c13 21 VSS 0.00271103f
r1 16 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.1195 $Y=0.2025 $X2=1.1320 $Y2=0.2025
r2 45 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.1170 $Y=0.2025 $X2=1.1195 $Y2=0.2025
r3 43 41 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0430 $Y=0.2025 $X2=1.0405 $Y2=0.2025
r4 2 41 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0260 $Y=0.2025 $X2=1.0405 $Y2=0.2025
r5 15 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0115 $Y=0.2025 $X2=1.0260 $Y2=0.2025
r6 42 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0090 $Y=0.2025 $X2=1.0115 $Y2=0.2025
r7 4 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.1340 $Y=0.2025
+ $X2=1.1340 $Y2=0.2340
r8 2 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0260 $Y=0.2025
+ $X2=1.0260 $Y2=0.2340
r9 38 39 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.1340
+ $Y=0.2340 $X2=1.1480 $Y2=0.2340
r10 37 38 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.0800
+ $Y=0.2340 $X2=1.1340 $Y2=0.2340
r11 36 37 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.2340 $X2=1.0800 $Y2=0.2340
r12 18 36 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.0145
+ $Y=0.2340 $X2=1.0260 $Y2=0.2340
r13 21 33 7.2121 $w=1.53211e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1620 $Y=0.2340 $X2=1.1620 $Y2=0.1960
r14 21 39 1.61554 $w=1.62143e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1620 $Y=0.2340 $X2=1.1480 $Y2=0.2340
r15 14 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.1195 $Y=0.0675 $X2=1.1320 $Y2=0.0675
r16 35 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.1170 $Y=0.0675 $X2=1.1195 $Y2=0.0675
r17 32 33 8.80291 $w=1.3e-08 $l=3.78e-08 $layer=M1 $thickness=3.6e-08 $X=1.1620
+ $Y=0.1582 $X2=1.1620 $Y2=0.1960
r18 31 32 2.15701 $w=1.3e-08 $l=9.2e-09 $layer=M1 $thickness=3.6e-08 $X=1.1620
+ $Y=0.1490 $X2=1.1620 $Y2=0.1582
r19 31 30 3.20636 $w=1.3e-08 $l=1.38e-08 $layer=M1 $thickness=3.6e-08 $X=1.1620
+ $Y=0.1490 $X2=1.1620 $Y2=0.1352
r20 19 20 9.4274 $w=1.48568e-08 $l=4.75e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1620 $Y=0.0835 $X2=1.1620 $Y2=0.0360
r21 19 30 12.0676 $w=1.3e-08 $l=5.17e-08 $layer=M1 $thickness=3.6e-08 $X=1.1620
+ $Y=0.0835 $X2=1.1620 $Y2=0.1352
r22 3 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.1340 $Y=0.0675
+ $X2=1.1340 $Y2=0.0360
r23 20 29 1.61554 $w=1.62143e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1620 $Y=0.0360 $X2=1.1480 $Y2=0.0360
r24 28 29 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.1340
+ $Y=0.0360 $X2=1.1480 $Y2=0.0360
r25 27 28 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.0800
+ $Y=0.0360 $X2=1.1340 $Y2=0.0360
r26 26 27 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.0360 $X2=1.0800 $Y2=0.0360
r27 17 26 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.0145
+ $Y=0.0360 $X2=1.0260 $Y2=0.0360
r28 1 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0260 $Y=0.0675
+ $X2=1.0260 $Y2=0.0360
r29 25 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.0430 $Y=0.0675 $X2=1.0405 $Y2=0.0675
r30 1 23 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.0260 $Y=0.0675 $X2=1.0405 $Y2=0.0675
r31 13 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.0115 $Y=0.0675 $X2=1.0260 $Y2=0.0675
r32 24 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.0090 $Y=0.0675 $X2=1.0115 $Y2=0.0675
.ends

.subckt PM_DFFHQNx3_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.00425975f
.ends

.subckt PM_DFFHQNx3_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.00416044f
.ends

.subckt PM_DFFHQNx3_ASAP7_75t_R%PD1 VSS 7 10 5 4 1
c1 1 VSS 0.0106264f
c2 4 VSS 0.00318963f
c3 5 VSS 0.00185363f
r1 10 9 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r2 8 9 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r3 5 8 0.123457 $w=8.1e-08 $l=1e-08 $layer=N_src_drn $thickness=1e-09 $X=0.3780
+ $Y=0.0675 $X2=0.3880 $Y2=0.0675
r4 4 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3220 $Y2=0.0675
r5 7 4 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r6 1 5 1e-05
.ends

.subckt PM_DFFHQNx3_ASAP7_75t_R%CLK VSS 10 3 8 5 1 6 7 4
c1 1 VSS 0.00247693f
c2 3 VSS 0.0596806f
c3 4 VSS 0.000948655f
c4 5 VSS 0.00400146f
c5 6 VSS 0.00388539f
c6 7 VSS 0.00220062f
c7 8 VSS 0.0020721f
r1 6 18 3.22357 $w=2.26279e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.2125 $X2=0.1080 $Y2=0.1820
r2 5 16 3.22357 $w=2.26279e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0575 $X2=0.1080 $Y2=0.0880
r3 17 18 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.1820 $X2=0.1080 $Y2=0.1820
r4 8 14 0.54189 $w=3.37e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1820 $X2=0.0810 $Y2=0.1630
r5 8 17 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1820 $X2=0.0945 $Y2=0.1820
r6 15 16 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.0880 $X2=0.1080 $Y2=0.0880
r7 7 15 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0880 $X2=0.0945 $Y2=0.0880
r8 13 14 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1530 $X2=0.0810 $Y2=0.1630
r9 12 13 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1530
r10 11 12 2.85657 $w=1.3e-08 $l=1.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1227 $X2=0.0810 $Y2=0.1350
r11 10 11 0.874462 $w=1.3e-08 $l=3.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1227
r12 10 4 1.57403 $w=1.3e-08 $l=6.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1122
r13 4 7 1.76614 $w=2.65738e-08 $l=2.42e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1122 $X2=0.0810 $Y2=0.0880
r14 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r15 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_DFFHQNx3_ASAP7_75t_R%D VSS 19 3 5 6 7 9 1 4 8
c1 1 VSS 0.0107701f
c2 3 VSS 0.0836248f
c3 4 VSS 0.00376895f
c4 5 VSS 0.00342498f
c5 6 VSS 0.00164304f
c6 7 VSS 0.00748512f
c7 8 VSS 0.00111109f
c8 9 VSS 0.00732006f
r1 9 21 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2430 $Y2=0.2140
r2 7 18 5.17411 $w=1.46514e-08 $l=2.72e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0360 $X2=0.2430 $Y2=0.0632
r3 5 8 7.7975 $w=1.41688e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1735 $X2=0.2430 $Y2=0.1350
r4 5 21 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1735 $X2=0.2430 $Y2=0.2140
r5 19 20 2.85657 $w=1.3e-08 $l=1.22e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0820 $X2=0.2430 $Y2=0.0942
r6 19 18 4.37231 $w=1.3e-08 $l=1.88e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0820 $X2=0.2430 $Y2=0.0632
r7 4 8 3.2503 $w=1.53684e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1160 $X2=0.2430 $Y2=0.1350
r8 4 20 5.07188 $w=1.3e-08 $l=2.18e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1160 $X2=0.2430 $Y2=0.0942
r9 16 17 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2715
+ $Y=0.1350 $X2=0.2810 $Y2=0.1350
r10 6 16 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2615
+ $Y=0.1350 $X2=0.2715 $Y2=0.1350
r11 6 8 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2615 $Y=0.1350 $X2=0.2430 $Y2=0.1350
r12 14 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2770 $Y=0.1350
+ $X2=0.2810 $Y2=0.1350
r13 12 14 4.43042 $w=1.53e-08 $l=7.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.2845 $Y=0.1350 $X2=0.2770 $Y2=0.1350
r14 1 11 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.2885
+ $Y=0.1350 $X2=0.2985 $Y2=0.1350
r15 1 12 1.86855 $w=1.78125e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.2885 $Y=0.1350 $X2=0.2845 $Y2=0.1350
r16 3 11 2.53453 $w=1.32811e-07 $l=1.5e-09 $layer=LIG $thickness=5.23243e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2985 $Y2=0.1350
r17 3 12 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2845 $Y2=0.1350
.ends

.subckt PM_DFFHQNx3_ASAP7_75t_R%PD3 VSS 2 4 1
c1 1 VSS 0.000972121f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0405 $X2=0.4905 $Y2=0.0405
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0405 $X2=0.4735 $Y2=0.0405
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4735 $Y=0.0405 $X2=0.4905 $Y2=0.0405
.ends

.subckt PM_DFFHQNx3_ASAP7_75t_R%PD4 VSS 2 4 1
c1 1 VSS 0.000945814f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.2295 $X2=0.7605 $Y2=0.2295
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.2295 $X2=0.7435 $Y2=0.2295
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7435 $Y=0.2295 $X2=0.7605 $Y2=0.2295
.ends

.subckt PM_DFFHQNx3_ASAP7_75t_R%PD5 VSS 7 12 4 1 5
c1 1 VSS 0.00741156f
c2 4 VSS 0.00187901f
c3 5 VSS 0.00237517f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.0405 $X2=0.7705 $Y2=0.0405
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7580 $Y=0.0405 $X2=0.7705 $Y2=0.0405
r3 9 5 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.7425
+ $Y=0.0405 $X2=0.7560 $Y2=0.0405
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.7275
+ $Y=0.0405 $X2=0.7425 $Y2=0.0405
r5 1 8 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.7020
+ $Y=0.0405 $X2=0.7275 $Y2=0.0405
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.0405 $X2=0.7000 $Y2=0.0405
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.0405 $X2=0.6875 $Y2=0.0405
.ends

.subckt PM_DFFHQNx3_ASAP7_75t_R%MH VSS 9 49 53 59 63 10 18 14 12 3 15 4 16 19
+ 17 20 1
c1 1 VSS 0.000361495f
c2 3 VSS 0.00584127f
c3 4 VSS 0.00560549f
c4 9 VSS 0.0363931f
c5 10 VSS 0.00226919f
c6 11 VSS 9.01132e-20
c7 12 VSS 0.00280436f
c8 13 VSS 6.90288e-20
c9 14 VSS 0.00883632f
c10 15 VSS 0.0013864f
c11 16 VSS 0.000721375f
c12 17 VSS 0.000427611f
c13 18 VSS 0.0060776f
c14 19 VSS 1.21202e-20
c15 20 VSS 0.00240131f
r1 63 62 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r2 61 62 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r3 3 61 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3760 $Y=0.2295 $X2=0.3880 $Y2=0.2295
r4 13 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2295 $X2=0.3760 $Y2=0.2295
r5 57 58 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r6 59 57 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.1890 $X2=0.3635 $Y2=0.1890
r7 12 58 0.185185 $w=5.4e-08 $l=1e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r8 12 3 0.518519 $w=3.9e-08 $l=4.05494e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.1890 $X2=0.3760 $Y2=0.2295
r9 3 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2295
+ $X2=0.3780 $Y2=0.2340
r10 53 52 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r11 51 52 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4420 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r12 4 51 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4300 $Y=0.0405 $X2=0.4420 $Y2=0.0405
r13 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0405 $X2=0.4300 $Y2=0.0405
r14 10 4 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0810 $X2=0.4300 $Y2=0.0810
r15 49 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0810 $X2=0.4175 $Y2=0.0810
r16 45 46 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r17 43 46 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r18 42 43 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4160
+ $Y=0.2340 $X2=0.4050 $Y2=0.2340
r19 14 20 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4340
+ $Y=0.2340 $X2=0.4590 $Y2=0.2340
r20 14 42 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4340
+ $Y=0.2340 $X2=0.4160 $Y2=0.2340
r21 4 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0405
+ $X2=0.4320 $Y2=0.0360
r22 20 34 3.01468 $w=1.741e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4590 $Y2=0.2140
r23 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4455 $Y2=0.0360
r24 18 31 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4590 $Y2=0.0630
r25 18 37 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4455 $Y2=0.0360
r26 33 34 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1850 $X2=0.4590 $Y2=0.2140
r27 32 33 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1660 $X2=0.4590 $Y2=0.1850
r28 16 19 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1525 $X2=0.4590 $Y2=0.1310
r29 16 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1525 $X2=0.4590 $Y2=0.1660
r30 30 31 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0900 $X2=0.4590 $Y2=0.0630
r31 29 30 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1025 $X2=0.4590 $Y2=0.0900
r32 15 19 2.78392 $w=1.56471e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1140 $X2=0.4590 $Y2=0.1310
r33 15 29 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1140 $X2=0.4590 $Y2=0.1025
r34 19 28 4.18306 $w=1.49565e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1310 $X2=0.4820 $Y2=0.1310
r35 27 28 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5000
+ $Y=0.1310 $X2=0.4820 $Y2=0.1310
r36 26 27 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1310 $X2=0.5000 $Y2=0.1310
r37 17 25 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1310 $X2=0.5670 $Y2=0.1310
r38 17 26 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1310 $X2=0.5130 $Y2=0.1310
r39 1 22 2.36633 $w=2.3e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.5670
+ $Y=0.1305 $X2=0.5670 $Y2=0.1305
r40 1 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1305
+ $X2=0.5670 $Y2=0.1310
r41 9 22 0.314665 $w=2.27e-07 $l=4.5e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5670 $Y=0.1350 $X2=0.5670 $Y2=0.1305
r42 3 12 1e-05
.ends

.subckt PM_DFFHQNx3_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.00485236f
.ends

.subckt PM_DFFHQNx3_ASAP7_75t_R%PU1 VSS 2 4 1
c1 1 VSS 0.000985137f
r1 4 3 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3365 $Y2=0.2025
r2 2 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3195 $Y2=0.2025
r3 1 3 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3195 $Y=0.2025 $X2=0.3365 $Y2=0.2025
.ends

.subckt PM_DFFHQNx3_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.00486835f
.ends

.subckt PM_DFFHQNx3_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.0415632f
.ends

.subckt PM_DFFHQNx3_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.0415747f
.ends

.subckt PM_DFFHQNx3_ASAP7_75t_R%PD2 VSS 7 12 4 5 1
c1 1 VSS 0.00730034f
c2 4 VSS 0.0018873f
c3 5 VSS 0.0023344f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4880 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r3 9 5 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.4605
+ $Y=0.2295 $X2=0.4860 $Y2=0.2295
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.4455
+ $Y=0.2295 $X2=0.4605 $Y2=0.2295
r5 1 8 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4320
+ $Y=0.2295 $X2=0.4455 $Y2=0.2295
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2295 $X2=0.4300 $Y2=0.2295
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2295 $X2=0.4175 $Y2=0.2295
.ends

.subckt PM_DFFHQNx3_ASAP7_75t_R%SS VSS 9 31 41 12 10 11 15 4 3 14 1 16 13
c1 1 VSS 0.00104865f
c2 3 VSS 0.00624362f
c3 4 VSS 0.00663132f
c4 9 VSS 0.0384418f
c5 10 VSS 0.00326636f
c6 11 VSS 0.00325094f
c7 12 VSS 0.00185094f
c8 13 VSS 0.0137729f
c9 14 VSS 0.00923421f
c10 15 VSS 0.00743183f
c11 16 VSS 0.0032393f
c12 17 VSS 0.00368061f
c13 18 VSS 0.00347458f
r1 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.2295 $X2=0.8620 $Y2=0.2295
r2 41 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.2295 $X2=0.8495 $Y2=0.2295
r3 4 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.2295
+ $X2=0.8640 $Y2=0.2340
r4 38 39 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.2340 $X2=0.8865 $Y2=0.2340
r5 14 18 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9180 $Y=0.2340 $X2=0.9450 $Y2=0.2340
r6 14 39 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.2340 $X2=0.8865 $Y2=0.2340
r7 18 36 0.56619 $w=2.22842e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.2340 $X2=0.9450 $Y2=0.2245
r8 35 36 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1975 $X2=0.9450 $Y2=0.2245
r9 34 35 6.64591 $w=1.3e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1690 $X2=0.9450 $Y2=0.1975
r10 33 34 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1445 $X2=0.9450 $Y2=0.1690
r11 32 33 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1195 $X2=0.9450 $Y2=0.1445
r12 15 17 8.84443 $w=1.496e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.0810 $X2=0.9450 $Y2=0.0360
r13 15 32 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.0810 $X2=0.9450 $Y2=0.1195
r14 10 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.0405 $X2=0.8620 $Y2=0.0405
r15 31 10 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.0405 $X2=0.8495 $Y2=0.0405
r16 17 29 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.0360 $X2=0.9180 $Y2=0.0360
r17 3 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.0405
+ $X2=0.8640 $Y2=0.0360
r18 28 29 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.0360 $X2=0.9180 $Y2=0.0360
r19 27 28 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.0360 $X2=0.8910 $Y2=0.0360
r20 26 27 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.0360 $X2=0.8640 $Y2=0.0360
r21 13 16 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.0360 $X2=0.7830 $Y2=0.0360
r22 13 26 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0360 $X2=0.8370 $Y2=0.0360
r23 12 23 8.04505 $w=1.3e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.0705 $X2=0.7830 $Y2=0.1050
r24 12 16 6.39593 $w=1.55565e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7830 $Y=0.0705 $X2=0.7830 $Y2=0.0360
r25 1 20 2.36633 $w=2.3e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.7830
+ $Y=0.1055 $X2=0.7830 $Y2=0.1055
r26 1 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7830 $Y=0.1055
+ $X2=0.7830 $Y2=0.1050
r27 9 20 0.314665 $w=2.27e-07 $l=2.95e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.7830 $Y=0.1350 $X2=0.7830 $Y2=0.1055
.ends

.subckt PM_DFFHQNx3_ASAP7_75t_R%MS VSS 10 41 44 48 50 13 17 18 14 3 15 12 1 11
+ 4 16
c1 1 VSS 0.00215636f
c2 3 VSS 0.0056759f
c3 4 VSS 0.00936263f
c4 10 VSS 0.037516f
c5 11 VSS 0.00302784f
c6 12 VSS 0.0028433f
c7 13 VSS 0.00240936f
c8 14 VSS 0.00185403f
c9 15 VSS 0.00401421f
c10 16 VSS 0.00177855f
c11 17 VSS 0.00124536f
c12 18 VSS 0.000447775f
c13 19 VSS 0.00278306f
r1 50 49 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.2295 $X2=0.6625 $Y2=0.2295
r2 13 49 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6500 $Y=0.2295 $X2=0.6625 $Y2=0.2295
r3 12 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2295 $X2=0.5920 $Y2=0.2295
r4 48 12 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.2295 $X2=0.5795 $Y2=0.2295
r5 45 13 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6210 $Y=0.2295 $X2=0.6480 $Y2=0.2295
r6 4 45 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08 $X=0.5940
+ $Y=0.2295 $X2=0.6210 $Y2=0.2295
r7 4 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2295
+ $X2=0.5940 $Y2=0.2340
r8 15 19 5.06479 $w=1.46038e-08 $l=2.70046e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5940 $Y=0.2340 $X2=0.6210 $Y2=0.2335
r9 44 43 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.0405 $X2=0.6085 $Y2=0.0405
r10 42 43 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6040 $Y=0.0405 $X2=0.6085 $Y2=0.0405
r11 3 42 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5920 $Y=0.0405 $X2=0.6040 $Y2=0.0405
r12 11 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.0405 $X2=0.5920 $Y2=0.0405
r13 41 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0405 $X2=0.5795 $Y2=0.0405
r14 19 36 0.983973 $w=1.77222e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.2335 $X2=0.6210 $Y2=0.2245
r15 3 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0405
+ $X2=0.5940 $Y2=0.0540
r16 35 36 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.2135 $X2=0.6210 $Y2=0.2245
r17 34 35 6.64591 $w=1.3e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1850 $X2=0.6210 $Y2=0.2135
r18 33 34 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1660 $X2=0.6210 $Y2=0.1850
r19 32 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1525 $X2=0.6210 $Y2=0.1660
r20 31 32 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1310 $X2=0.6210 $Y2=0.1525
r21 30 31 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1115 $X2=0.6210 $Y2=0.1310
r22 17 28 1.15159 $w=1.75e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1000 $X2=0.6210 $Y2=0.0900
r23 17 30 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1000 $X2=0.6210 $Y2=0.1115
r24 16 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0540 $X2=0.5940 $Y2=0.0720
r25 27 28 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6075 $Y=0.0900 $X2=0.6210 $Y2=0.0900
r26 18 26 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5940 $Y=0.0900 $X2=0.5805 $Y2=0.0900
r27 18 27 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5940 $Y=0.0900 $X2=0.6075 $Y2=0.0900
r28 18 29 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0900 $X2=0.5940 $Y2=0.0720
r29 25 26 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5490
+ $Y=0.0900 $X2=0.5805 $Y2=0.0900
r30 24 25 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0900 $X2=0.5490 $Y2=0.0900
r31 14 24 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5000
+ $Y=0.0900 $X2=0.5130 $Y2=0.0900
r32 1 21 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.5130
+ $Y=0.0900 $X2=0.5130 $Y2=0.0900
r33 1 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.0900
+ $X2=0.5130 $Y2=0.0900
r34 10 21 0.314665 $w=2.27e-07 $l=4.5e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5130 $Y2=0.0900
.ends

.subckt PM_DFFHQNx3_ASAP7_75t_R%CLKB VSS 14 15 16 17 81 83 18 20 26 6 7 23 24 4
+ 25 22 19 1 21 8 2
c1 1 VSS 0.00176254f
c2 2 VSS 0.000788121f
c3 3 VSS 0.000739371f
c4 4 VSS 0.00113479f
c5 6 VSS 0.00882486f
c6 7 VSS 0.00854139f
c7 8 VSS 0.00501353f
c8 14 VSS 0.00604138f
c9 15 VSS 0.00579999f
c10 16 VSS 0.00508597f
c11 17 VSS 0.00591633f
c12 18 VSS 0.00543717f
c13 19 VSS 0.00543076f
c14 20 VSS 0.00408362f
c15 21 VSS 0.00332498f
c16 22 VSS 0.00280899f
c17 23 VSS 0.00685649f
c18 24 VSS 0.00606705f
c19 25 VSS 0.0012541f
c20 26 VSS 0.00548571f
r1 19 7 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1600 $Y2=0.2160
r2 83 19 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r3 18 6 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1600 $Y2=0.0540
r4 81 18 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r5 4 79 2.78395 $w=2.4e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08 $X=0.7290
+ $Y=0.1780 $X2=0.7250 $Y2=0.1780
r6 17 4 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.7290 $Y=0.1350 $X2=0.7290 $Y2=0.1780
r7 3 72 10.3807 $w=2.30357e-08 $l=0 $layer=LISD $thickness=3.675e-08 $X=0.6210
+ $Y=0.1780 $X2=0.6210 $Y2=0.1780
r8 16 3 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.6210 $Y=0.1350 $X2=0.6210 $Y2=0.1780
r9 2 65 2.78395 $w=2.4e-08 $l=5e-09 $layer=LIG $thickness=4.8e-08 $X=0.4590
+ $Y=0.1780 $X2=0.4640 $Y2=0.1780
r10 15 2 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4590 $Y2=0.1780
r11 7 57 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1655 $Y2=0.2340
r12 6 53 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1655 $Y2=0.0360
r13 78 79 4.8113 $w=2.22e-08 $l=1.5e-09 $layer=LISD $thickness=2.7e-08
+ $X=0.7235 $Y=0.1780 $X2=0.7250 $Y2=0.1780
r14 77 78 10.8887 $w=2.22e-08 $l=2.15e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7020 $Y=0.1780 $X2=0.7235 $Y2=0.1780
r15 76 77 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6885 $Y=0.1780 $X2=0.7020 $Y2=0.1780
r16 75 76 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6750 $Y=0.1780 $X2=0.6885 $Y2=0.1780
r17 74 75 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6615 $Y=0.1780 $X2=0.6750 $Y2=0.1780
r18 73 74 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6480 $Y=0.1780 $X2=0.6615 $Y2=0.1780
r19 72 73 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6210 $Y=0.1780 $X2=0.6480 $Y2=0.1780
r20 71 72 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5940 $Y=0.1780 $X2=0.6210 $Y2=0.1780
r21 70 71 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5805 $Y=0.1780 $X2=0.5940 $Y2=0.1780
r22 69 70 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5670 $Y=0.1780 $X2=0.5805 $Y2=0.1780
r23 68 69 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5535 $Y=0.1780 $X2=0.5670 $Y2=0.1780
r24 67 68 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5400 $Y=0.1780 $X2=0.5535 $Y2=0.1780
r25 66 67 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5265 $Y=0.1780 $X2=0.5400 $Y2=0.1780
r26 64 65 10.3823 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4775 $Y=0.1780 $X2=0.4640 $Y2=0.1780
r27 63 64 11.142 $w=2.22e-08 $l=2.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4995 $Y=0.1780 $X2=0.4775 $Y2=0.1780
r28 62 66 1.51936 $w=2.22e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.5235
+ $Y=0.1780 $X2=0.5265 $Y2=0.1780
r29 61 62 5.31775 $w=2.22e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5130 $Y=0.1780 $X2=0.5235 $Y2=0.1780
r30 8 61 5.31775 $w=2.22e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5025 $Y=0.1780 $X2=0.5130 $Y2=0.1780
r31 8 63 1.51936 $w=2.22e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.5025
+ $Y=0.1780 $X2=0.4995 $Y2=0.1780
r32 57 58 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1655
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r33 24 50 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2340 $X2=0.1890 $Y2=0.2125
r34 24 58 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2340 $X2=0.1755 $Y2=0.2340
r35 53 54 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1655
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r36 23 49 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1890 $Y2=0.0575
r37 23 54 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1755 $Y2=0.0360
r38 51 61 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5130 $Y=0.1845
+ $X2=0.5130 $Y2=0.1780
r39 22 51 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1680 $X2=0.5130 $Y2=0.1845
r40 48 49 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0880 $X2=0.1890 $Y2=0.0575
r41 47 48 11.3097 $w=1.3e-08 $l=4.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1365 $X2=0.1890 $Y2=0.0880
r42 46 50 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1990 $X2=0.1890 $Y2=0.2125
r43 45 46 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1890 $X2=0.1890 $Y2=0.1990
r44 20 45 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1735 $X2=0.1890 $Y2=0.1890
r45 20 47 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1735 $X2=0.1890 $Y2=0.1365
r46 43 51 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.5130 $Y=0.1890
+ $X2=0.5130 $Y2=0.1845
r47 42 43 22.0364 $w=1.3e-08 $l=9.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.4185
+ $Y=0.1890 $X2=0.5130 $Y2=0.1890
r48 41 42 22.0364 $w=1.3e-08 $l=9.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1890 $X2=0.4185 $Y2=0.1890
r49 40 41 15.7403 $w=1.3e-08 $l=6.75e-08 $layer=M2 $thickness=3.6e-08 $X=0.2565
+ $Y=0.1890 $X2=0.3240 $Y2=0.1890
r50 39 40 15.7403 $w=1.3e-08 $l=6.75e-08 $layer=M2 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1890 $X2=0.2565 $Y2=0.1890
r51 39 45 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1890 $Y=0.1890
+ $X2=0.1890 $Y2=0.1890
r52 26 39 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.1775
+ $Y=0.1890 $X2=0.1890 $Y2=0.1890
r53 37 41 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.3240 $Y=0.1890
+ $X2=0.3240 $Y2=0.1890
r54 36 37 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1735 $X2=0.3240 $Y2=0.1890
r55 21 34 3.60008 $w=1.51951e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3240 $Y=0.1555 $X2=0.3240 $Y2=0.1350
r56 21 36 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1555 $X2=0.3240 $Y2=0.1735
r57 25 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r58 25 34 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3375 $Y=0.1350 $X2=0.3240 $Y2=0.1350
r59 14 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r60 1 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
.ends

.subckt PM_DFFHQNx3_ASAP7_75t_R%SH VSS 11 12 13 14 81 84 89 92 30 6 20 16 15 25
+ 27 18 19 17 5 23 29 2 28 24 22 1 26 21
c1 1 VSS 0.00260407f
c2 2 VSS 0.0154829f
c3 5 VSS 0.00683511f
c4 6 VSS 0.00674942f
c5 11 VSS 0.0383606f
c6 12 VSS 0.0821136f
c7 13 VSS 0.0813811f
c8 14 VSS 0.081091f
c9 15 VSS 0.00485332f
c10 16 VSS 0.00507605f
c11 17 VSS 0.00851979f
c12 18 VSS 0.00198004f
c13 19 VSS 0.00210104f
c14 20 VSS 0.00249636f
c15 21 VSS 0.00124119f
c16 22 VSS 0.00135985f
c17 23 VSS 0.00244906f
c18 24 VSS 0.0034666f
c19 25 VSS 0.00655629f
c20 26 VSS 0.00318495f
c21 27 VSS 0.00100235f
c22 28 VSS 0.00121936f
c23 29 VSS 0.00115755f
c24 30 VSS 0.00350322f
r1 92 91 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r2 5 91 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6500 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r3 88 5 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6380 $Y=0.0405 $X2=0.6500 $Y2=0.0405
r4 15 88 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0405 $X2=0.6380 $Y2=0.0405
r5 89 15 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.0405 $X2=0.6335 $Y2=0.0405
r6 14 75 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=1.1070
+ $Y=0.1350 $X2=1.1070 $Y2=0.1360
r7 13 69 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=1.0530
+ $Y=0.1350 $X2=1.0530 $Y2=0.1360
r8 12 61 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.9990 $Y=0.1350 $X2=0.9990 $Y2=0.1360
r9 84 83 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r10 82 83 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7120 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r11 6 82 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7000 $Y=0.2295 $X2=0.7120 $Y2=0.2295
r12 16 6 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.2295 $X2=0.7000 $Y2=0.2295
r13 81 16 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.2295 $X2=0.6875 $Y2=0.2295
r14 5 59 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.0405
+ $X2=0.6480 $Y2=0.0360
r15 73 75 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.0945 $Y=0.1360 $X2=1.1070 $Y2=0.1360
r16 72 73 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.0800 $Y=0.1360 $X2=1.0945 $Y2=0.1360
r17 70 72 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.0655 $Y=0.1360 $X2=1.0800 $Y2=0.1360
r18 69 70 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.0530 $Y=0.1360 $X2=1.0655 $Y2=0.1360
r19 67 69 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.0405 $Y=0.1360 $X2=1.0530 $Y2=0.1360
r20 66 67 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.0260 $Y=0.1360 $X2=1.0405 $Y2=0.1360
r21 64 66 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.0115 $Y=0.1360 $X2=1.0260 $Y2=0.1360
r22 62 64 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=1.0085 $Y=0.1360 $X2=1.0115 $Y2=0.1360
r23 61 62 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.9990
+ $Y=0.1360 $X2=1.0085 $Y2=0.1360
r24 2 61 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.9895
+ $Y=0.1360 $X2=0.9990 $Y2=0.1360
r25 6 52 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7020 $Y=0.2295
+ $X2=0.7020 $Y2=0.2330
r26 59 60 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6480
+ $Y=0.0360 $X2=0.6615 $Y2=0.0360
r27 57 60 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0360 $X2=0.6615 $Y2=0.0360
r28 56 57 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6860
+ $Y=0.0360 $X2=0.6750 $Y2=0.0360
r29 17 26 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.7040
+ $Y=0.0360 $X2=0.7290 $Y2=0.0360
r30 17 56 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7040
+ $Y=0.0360 $X2=0.6860 $Y2=0.0360
r31 54 61 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.9990 $Y=0.1445
+ $X2=0.9990 $Y2=0.1360
r32 24 54 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.9990
+ $Y=0.1245 $X2=0.9990 $Y2=0.1445
r33 52 53 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.2330 $X2=0.7155 $Y2=0.2330
r34 25 53 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.2330 $X2=0.7155 $Y2=0.2330
r35 26 45 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.0360 $X2=0.7290 $Y2=0.0630
r36 49 54 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.9990 $Y=0.1530
+ $X2=0.9990 $Y2=0.1445
r37 48 49 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1530 $X2=0.9990 $Y2=0.1530
r38 47 48 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1530 $X2=0.9450 $Y2=0.1530
r39 30 47 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.8795
+ $Y=0.1530 $X2=0.8910 $Y2=0.1530
r40 46 47 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.8910 $Y=0.1485 $X2=0.8910
+ $Y2=0.1530
r41 23 46 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1305 $X2=0.8910 $Y2=0.1485
r42 19 40 6.38362 $w=1.33509e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1975 $X2=0.7290 $Y2=0.1690
r43 19 25 7.09793 $w=1.42676e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1975 $X2=0.7290 $Y2=0.2330
r44 44 45 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.0900 $X2=0.7290 $Y2=0.0630
r45 43 44 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1000 $X2=0.7290 $Y2=0.0900
r46 42 43 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1100 $X2=0.7290 $Y2=0.1000
r47 18 27 4.67854 $w=1.44583e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1360 $X2=0.7290 $Y2=0.1600
r48 18 42 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1360 $X2=0.7290 $Y2=0.1100
r49 29 41 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1575 $X2=0.8910 $Y2=0.1665
r50 29 46 1.50855 $w=1.55e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1575 $X2=0.8910 $Y2=0.1485
r51 29 47 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.8910 $Y=0.1575 $X2=0.8910
+ $Y2=0.1530
r52 27 40 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1600 $X2=0.7290 $Y2=0.1690
r53 39 41 4.19024 $w=1.156e-08 $l=2.54018e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8660 $Y=0.1620 $X2=0.8910 $Y2=0.1665
r54 22 28 1.38478 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8480 $Y=0.1620 $X2=0.8370 $Y2=0.1620
r55 22 39 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8480
+ $Y=0.1620 $X2=0.8660 $Y2=0.1620
r56 38 40 4.4015 $w=1.35e-08 $l=2.78927e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7560 $Y=0.1620 $X2=0.7290 $Y2=0.1690
r57 37 38 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1620 $X2=0.7560 $Y2=0.1620
r58 20 28 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.1620 $X2=0.8370 $Y2=0.1620
r59 20 37 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.1620 $X2=0.7830 $Y2=0.1620
r60 28 36 4.88263 $w=1.47308e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8370 $Y=0.1620 $X2=0.8370 $Y2=0.1360
r61 21 36 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1180 $X2=0.8370 $Y2=0.1360
r62 11 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.8370
+ $Y=0.1350 $X2=0.8370 $Y2=0.1350
r63 1 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8370 $Y=0.1350
+ $X2=0.8370 $Y2=0.1360
.ends

.subckt PM_DFFHQNx3_ASAP7_75t_R%CLKN VSS 13 14 15 77 79 22 8 26 7 16 17 1 19 21
+ 20 18 28 23 2 24 3
c1 1 VSS 0.001618f
c2 2 VSS 4.49461e-20
c3 3 VSS 0.000195395f
c4 7 VSS 0.00749348f
c5 8 VSS 0.00762177f
c6 13 VSS 0.0596117f
c7 14 VSS 0.00439493f
c8 15 VSS 0.0045813f
c9 16 VSS 0.00603668f
c10 17 VSS 0.00596318f
c11 18 VSS 0.00537565f
c12 19 VSS 0.0035035f
c13 20 VSS 0.00462689f
c14 21 VSS 0.00451543f
c15 22 VSS 0.000592632f
c16 23 VSS 0.000586274f
c17 24 VSS 0.00132874f
c18 25 VSS 0.00366894f
c19 26 VSS 0.00155567f
c20 27 VSS 0.00379262f
c21 28 VSS 0.0239016f
r1 79 78 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r2 17 78 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r3 77 76 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r4 16 76 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r5 8 74 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0550 $Y2=0.2340
r6 7 71 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0550 $Y2=0.0360
r7 73 74 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.2340 $X2=0.0550 $Y2=0.2340
r8 21 73 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0460 $Y2=0.2340
r9 21 27 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0180 $Y2=0.2340
r10 70 71 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.0360 $X2=0.0550 $Y2=0.0360
r11 20 70 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0460 $Y2=0.0360
r12 20 25 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0180 $Y2=0.0360
r13 27 63 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.2340 $X2=0.0180 $Y2=0.2125
r14 25 61 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.0360 $X2=0.0180 $Y2=0.0575
r15 3 58 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6750 $Y=0.1350
+ $X2=0.6750 $Y2=0.1440
r16 15 3 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6750
+ $Y=0.1350 $X2=0.6750 $Y2=0.1350
r17 2 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
r18 14 2 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r19 62 63 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1820 $X2=0.0180 $Y2=0.2125
r20 19 26 0.998523 $w=1.74118e-08 $l=1.01119e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1630 $X2=0.0165 $Y2=0.1530
r21 19 62 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1630 $X2=0.0180 $Y2=0.1820
r22 60 61 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0880 $X2=0.0180 $Y2=0.0575
r23 18 26 5.19594 $w=1.44151e-08 $l=2.80401e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1250 $X2=0.0165 $Y2=0.1530
r24 18 60 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1250 $X2=0.0180 $Y2=0.0880
r25 24 58 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1135 $X2=0.6750 $Y2=0.1440
r26 23 56 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1530
r27 52 53 1.90199 $w=1.38333e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.0255 $Y=0.1530 $X2=0.0345 $Y2=0.1530
r28 26 52 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0165
+ $Y=0.1530 $X2=0.0255 $Y2=0.1530
r29 50 58 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.6750 $Y=0.1530
+ $X2=0.6750 $Y2=0.1440
r30 49 50 18.3054 $w=1.3e-08 $l=7.85e-08 $layer=M2 $thickness=3.6e-08 $X=0.5965
+ $Y=0.1530 $X2=0.6750 $Y2=0.1530
r31 48 49 29.3819 $w=1.3e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.4705
+ $Y=0.1530 $X2=0.5965 $Y2=0.1530
r32 47 48 15.2739 $w=1.3e-08 $l=6.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1530 $X2=0.4705 $Y2=0.1530
r33 47 56 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4050 $Y=0.1530
+ $X2=0.4050 $Y2=0.1530
r34 46 47 27.8662 $w=1.3e-08 $l=1.195e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.2855 $Y=0.1530 $X2=0.4050 $Y2=0.1530
r35 45 46 27.5164 $w=1.3e-08 $l=1.18e-07 $layer=M2 $thickness=3.6e-08 $X=0.1675
+ $Y=0.1530 $X2=0.2855 $Y2=0.1530
r36 44 45 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M2 $thickness=3.6e-08 $X=0.1510
+ $Y=0.1530 $X2=0.1675 $Y2=0.1530
r37 43 44 13.7582 $w=1.3e-08 $l=5.9e-08 $layer=M2 $thickness=3.6e-08 $X=0.0920
+ $Y=0.1530 $X2=0.1510 $Y2=0.1530
r38 42 43 13.7582 $w=1.3e-08 $l=5.9e-08 $layer=M2 $thickness=3.6e-08 $X=0.0330
+ $Y=0.1530 $X2=0.0920 $Y2=0.1530
r39 42 53 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.0330 $Y=0.1530
+ $X2=0.0345 $Y2=0.1530
r40 28 42 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.0215
+ $Y=0.1530 $X2=0.0330 $Y2=0.1530
r41 39 44 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1510 $Y=0.1440
+ $X2=0.1510 $Y2=0.1530
r42 22 39 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1510
+ $Y=0.1160 $X2=0.1510 $Y2=0.1440
r43 37 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1550 $Y=0.1350
+ $X2=0.1510 $Y2=0.1440
r44 36 37 4.43042 $w=1.53e-08 $l=7.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1475 $Y=0.1350 $X2=0.1550 $Y2=0.1350
r45 34 36 1.86855 $w=1.78125e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1435 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r46 1 34 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.1335
+ $Y=0.1350 $X2=0.1435 $Y2=0.1350
r47 13 1 2.53453 $w=1.32811e-07 $l=1.5e-09 $layer=LIG $thickness=5.23243e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1335 $Y2=0.1350
r48 13 36 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r49 8 17 1e-05
r50 7 16 1e-05
.ends


*
.SUBCKT DFFHQNx3_ASAP7_75t_R VSS VDD CLK D QN
*
* VSS VSS
* VDD VDD
* CLK CLK
* D D
* QN QN
*
*

MM20 N_MM20_d N_MM20_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM23 N_MM23_d N_MM22_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM10_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM6 N_MM6_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM12 N_MM12_d N_MM12_g N_MM12_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM17 N_MM17_d N_MM13_g N_MM17_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM16 N_MM16_d N_MM19_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM14 N_MM14_d N_MM14_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM24 N_MM24_d N_MM24_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@3 N_MM24@3_d N_MM24@3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@2 N_MM24@2_d N_MM24@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM21 N_MM21_d N_MM20_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM22 N_MM22_d N_MM22_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM13 N_MM13_d N_MM13_g N_MM13_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM18 N_MM18_d N_MM18_g N_MM18_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM19 N_MM19_d N_MM19_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM15 N_MM15_d N_MM14_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM25 N_MM25_d N_MM24_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@3 N_MM25@3_d N_MM24@3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@2 N_MM25@2_d N_MM24@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "DFFHQNx3_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "DFFHQNx3_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_DFFHQNx3_ASAP7_75t_R%noxref_27 VSS N_noxref_27_1
+ PM_DFFHQNx3_ASAP7_75t_R%noxref_27
cc_1 N_noxref_27_1 N_SS_11 0.000639303f
cc_2 N_noxref_27_1 N_MM24_g 0.00172026f
cc_3 N_noxref_27_1 N_noxref_24_1 0.000477825f
cc_4 N_noxref_27_1 N_noxref_25_1 0.00776243f
cc_5 N_noxref_27_1 N_noxref_26_1 0.00123288f
x_PM_DFFHQNx3_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_DFFHQNx3_ASAP7_75t_R%noxref_24
cc_6 N_noxref_24_1 N_SS_10 0.0170327f
cc_7 N_noxref_24_1 N_SH_1 0.000196229f
cc_8 N_noxref_24_1 N_MM14_g 0.00593676f
x_PM_DFFHQNx3_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_DFFHQNx3_ASAP7_75t_R%noxref_25
cc_9 N_noxref_25_1 N_SS_11 0.0169151f
cc_10 N_noxref_25_1 N_SH_1 0.000200836f
cc_11 N_noxref_25_1 N_MM14_g 0.00603601f
cc_12 N_noxref_25_1 N_noxref_24_1 0.0015414f
x_PM_DFFHQNx3_ASAP7_75t_R%noxref_29 VSS N_noxref_29_1
+ PM_DFFHQNx3_ASAP7_75t_R%noxref_29
cc_13 N_noxref_29_1 N_MM24@2_g 0.00147713f
cc_14 N_noxref_29_1 N_QN_16 0.0378708f
cc_15 N_noxref_29_1 N_noxref_28_1 0.00176784f
x_PM_DFFHQNx3_ASAP7_75t_R%noxref_28 VSS N_noxref_28_1
+ PM_DFFHQNx3_ASAP7_75t_R%noxref_28
cc_16 N_noxref_28_1 N_MM24@2_g 0.00147623f
cc_17 N_noxref_28_1 N_QN_14 0.037595f
x_PM_DFFHQNx3_ASAP7_75t_R%noxref_26 VSS N_noxref_26_1
+ PM_DFFHQNx3_ASAP7_75t_R%noxref_26
cc_18 N_noxref_26_1 N_SS_10 0.000658809f
cc_19 N_noxref_26_1 N_MM24_g 0.0017013f
cc_20 N_noxref_26_1 N_noxref_24_1 0.00776096f
cc_21 N_noxref_26_1 N_noxref_25_1 0.000476381f
x_PM_DFFHQNx3_ASAP7_75t_R%QN VSS QN N_MM24_d N_MM24@3_d N_MM24@2_d N_MM25_d
+ N_MM25@3_d N_MM25@2_d N_QN_13 N_QN_19 N_QN_18 N_QN_15 N_QN_3 N_QN_4 N_QN_2
+ N_QN_1 N_QN_16 N_QN_14 PM_DFFHQNx3_ASAP7_75t_R%QN
cc_22 N_QN_13 N_SH_24 0.000229275f
cc_23 N_QN_13 N_MM24@2_g 0.00148455f
cc_24 N_QN_13 N_SH_2 0.000469939f
cc_25 N_QN_13 N_SH_30 0.000725327f
cc_26 N_QN_19 N_SH_2 0.00077582f
cc_27 N_QN_18 N_MM24@2_g 0.000812562f
cc_28 N_QN_15 N_MM24@3_g 0.0308554f
cc_29 N_QN_3 N_MM24@2_g 0.000867566f
cc_30 N_QN_4 N_MM24@2_g 0.000904378f
cc_31 N_QN_2 N_SH_24 0.000907531f
cc_32 N_QN_1 N_MM24@3_g 0.00199954f
cc_33 N_QN_2 N_MM24@3_g 0.00214847f
cc_34 N_QN_16 N_MM24@2_g 0.0151504f
cc_35 N_QN_15 N_SH_2 0.00693895f
cc_36 N_QN_14 N_MM24@2_g 0.0524462f
cc_37 N_QN_13 N_MM24_g 0.0372032f
cc_38 N_QN_13 N_MM24@3_g 0.0684768f
x_PM_DFFHQNx3_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_DFFHQNx3_ASAP7_75t_R%noxref_18
cc_39 N_noxref_18_1 N_MM20_g 0.0036837f
cc_40 N_noxref_18_1 N_CLKN_19 6.24368e-20
cc_41 N_noxref_18_1 N_CLKN_18 0.000315549f
cc_42 N_noxref_18_1 N_CLKN_7 0.000503374f
cc_43 N_noxref_18_1 N_CLKN_16 0.0278219f
x_PM_DFFHQNx3_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_DFFHQNx3_ASAP7_75t_R%noxref_19
cc_44 N_noxref_19_1 N_MM20_g 0.00367249f
cc_45 N_noxref_19_1 N_CLKN_26 8.87656e-20
cc_46 N_noxref_19_1 N_CLKN_18 0.000153431f
cc_47 N_noxref_19_1 N_CLKN_19 0.000196766f
cc_48 N_noxref_19_1 N_CLKN_8 0.000505002f
cc_49 N_noxref_19_1 N_CLKN_17 0.0278547f
cc_50 N_noxref_19_1 N_noxref_18_1 0.00204748f
x_PM_DFFHQNx3_ASAP7_75t_R%PD1 VSS N_MM5_d N_MM4_s N_PD1_5 N_PD1_4 N_PD1_1
+ PM_DFFHQNx3_ASAP7_75t_R%PD1
cc_51 N_PD1_5 N_CLKN_2 0.000858369f
cc_52 N_PD1_5 N_CLKN_23 0.000316652f
cc_53 N_PD1_5 N_MM10_g 0.0343289f
cc_54 N_PD1_4 N_MM3_g 0.0359294f
cc_55 N_PD1_5 N_CLKB_25 0.000413009f
cc_56 N_PD1_5 N_CLKB_1 0.00234471f
cc_57 N_PD1_5 N_MM1_g 0.0735623f
cc_58 N_PD1_1 N_MH_4 0.00122241f
cc_59 N_PD1_1 N_MH_10 0.00350019f
x_PM_DFFHQNx3_ASAP7_75t_R%CLK VSS CLK N_MM20_g N_CLK_8 N_CLK_5 N_CLK_1 N_CLK_6
+ N_CLK_7 N_CLK_4 PM_DFFHQNx3_ASAP7_75t_R%CLK
x_PM_DFFHQNx3_ASAP7_75t_R%D VSS D N_MM3_g N_D_5 N_D_6 N_D_7 N_D_9 N_D_1 N_D_4
+ N_D_8 PM_DFFHQNx3_ASAP7_75t_R%D
cc_60 N_D_5 N_CLKN_22 0.000146036f
cc_61 N_D_5 N_CLKN_23 7.47542e-20
cc_62 N_D_5 N_CLKN_1 0.000102901f
cc_63 N_D_6 N_CLKN_28 0.000655933f
cc_64 N_D_5 N_CLKN_28 0.00334804f
x_PM_DFFHQNx3_ASAP7_75t_R%PD3 VSS N_MM9_s N_MM8_d N_PD3_1
+ PM_DFFHQNx3_ASAP7_75t_R%PD3
cc_65 N_PD3_1 N_MM9_g 0.00773035f
cc_66 N_PD3_1 N_MM11_g 0.00773412f
x_PM_DFFHQNx3_ASAP7_75t_R%PD4 VSS N_MM18_s N_MM19_d N_PD4_1
+ PM_DFFHQNx3_ASAP7_75t_R%PD4
cc_67 N_PD4_1 N_MM18_g 0.00773066f
cc_68 N_PD4_1 N_MM19_g 0.00776505f
x_PM_DFFHQNx3_ASAP7_75t_R%PD5 VSS N_MM17_s N_MM16_d N_PD5_4 N_PD5_1 N_PD5_5
+ PM_DFFHQNx3_ASAP7_75t_R%PD5
cc_69 N_PD5_4 N_MM13_g 0.0152671f
cc_70 N_PD5_1 N_MM18_g 0.000759258f
cc_71 N_PD5_4 N_MM18_g 0.00694996f
cc_72 N_PD5_5 N_MM18_g 0.0239775f
cc_73 N_PD5_1 N_MM19_g 0.000915782f
cc_74 N_PD5_5 N_MM19_g 0.0155365f
cc_75 N_PD5_1 N_SH_15 0.000516159f
cc_76 N_PD5_1 N_SH_17 0.000448338f
cc_77 N_PD5_1 N_SH_18 0.000599439f
cc_78 N_PD5_4 N_SH_5 0.000664227f
cc_79 N_PD5_1 N_SH_26 0.00238643f
x_PM_DFFHQNx3_ASAP7_75t_R%MH VSS N_MM7_g N_MM4_d N_MM9_d N_MM1_d N_MM10_d
+ N_MH_10 N_MH_18 N_MH_14 N_MH_12 N_MH_3 N_MH_15 N_MH_4 N_MH_16 N_MH_19 N_MH_17
+ N_MH_20 N_MH_1 PM_DFFHQNx3_ASAP7_75t_R%MH
cc_80 N_MH_10 N_CLKN_3 0.000103934f
cc_81 N_MH_10 N_CLKN_28 0.000117104f
cc_82 N_MH_10 N_MM13_g 0.000188959f
cc_83 N_MH_10 N_CLKN_23 0.000326569f
cc_84 N_MH_18 N_CLKN_23 0.000369724f
cc_85 N_MH_14 N_CLKN_23 0.000396021f
cc_86 N_MH_12 N_MM10_g 0.016425f
cc_87 N_MH_3 N_CLKN_2 0.000773759f
cc_88 N_MH_15 N_CLKN_23 0.00110459f
cc_89 N_MH_4 N_MM10_g 0.00111959f
cc_90 N_MH_3 N_MM10_g 0.00123236f
cc_91 N_MH_16 N_CLKN_23 0.00124343f
cc_92 N_MH_10 N_CLKN_2 0.00164744f
cc_93 N_MH_19 N_CLKN_23 0.00296626f
cc_94 N_MH_17 N_CLKN_28 0.0035162f
cc_95 N_MH_10 N_MM10_g 0.0529684f
cc_96 N_MH_10 N_CLKB_22 0.000365996f
cc_97 N_MH_10 N_MM1_g 0.000402217f
cc_98 N_MH_10 N_CLKB_21 0.00017697f
cc_99 N_MH_10 N_CLKB_25 0.000272618f
cc_100 N_MH_20 N_CLKB_22 0.000316163f
cc_101 N_MH_16 N_CLKB_22 0.00266696f
cc_102 N_MH_3 N_CLKB_1 0.000337994f
cc_103 N_MH_17 N_CLKB_8 0.000557321f
cc_104 N_MH_4 N_MM9_g 0.000623503f
cc_105 N_MH_3 N_CLKB_21 0.000652426f
cc_106 N_MH_1 N_CLKB_8 0.00227377f
cc_107 N_MH_16 N_CLKB_2 0.000779248f
cc_108 N_MH_12 N_CLKB_1 0.000794579f
cc_109 N_MH_3 N_MM1_g 0.00175451f
cc_110 N_MH_14 N_CLKB_26 0.00280152f
cc_111 N_MH_17 N_CLKB_22 0.00357965f
cc_112 N_MM7_g N_CLKB_8 0.00464828f
cc_113 N_MH_12 N_MM1_g 0.033696f
cc_114 N_MM7_g N_MM12_g 0.0127424f
cc_115 N_MH_10 N_MM9_g 0.0364081f
cc_116 N_MH_17 N_MM11_g 0.000358875f
cc_117 N_MH_4 N_MS_1 0.000395717f
cc_118 N_MH_17 N_MS_1 0.000829706f
cc_119 N_MM7_g N_MS_3 0.000906615f
cc_120 N_MH_1 N_MS_14 0.000924777f
cc_121 N_MH_17 N_MS_17 0.00101626f
cc_122 N_MH_1 N_MM11_g 0.00114166f
cc_123 N_MM7_g N_MS_1 0.00116098f
cc_124 N_MH_15 N_MS_14 0.00124188f
cc_125 N_MM7_g N_MS_12 0.00639278f
cc_126 N_MM7_g N_MS_11 0.00641085f
cc_127 N_MH_17 N_MS_14 0.00738548f
cc_128 N_MM7_g N_MM11_g 0.0293738f
x_PM_DFFHQNx3_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_DFFHQNx3_ASAP7_75t_R%noxref_20
cc_129 N_noxref_20_1 N_CLKN_1 0.000398066f
cc_130 N_noxref_20_1 N_MM22_g 0.00343386f
cc_131 N_noxref_20_1 N_CLKB_6 0.000423111f
cc_132 N_noxref_20_1 N_CLKB_18 0.0270308f
x_PM_DFFHQNx3_ASAP7_75t_R%PU1 VSS N_MM3_d N_MM1_s N_PU1_1
+ PM_DFFHQNx3_ASAP7_75t_R%PU1
cc_133 N_PU1_1 N_MM3_g 0.0171044f
cc_134 N_PU1_1 N_MM1_g 0.0169733f
x_PM_DFFHQNx3_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_DFFHQNx3_ASAP7_75t_R%noxref_21
cc_135 N_noxref_21_1 N_CLKN_1 0.000396541f
cc_136 N_noxref_21_1 N_MM22_g 0.00344681f
cc_137 N_noxref_21_1 N_CLKB_7 0.000426471f
cc_138 N_noxref_21_1 N_CLKB_19 0.0270307f
cc_139 N_noxref_21_1 N_noxref_20_1 0.00141787f
x_PM_DFFHQNx3_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_DFFHQNx3_ASAP7_75t_R%noxref_22
cc_140 N_noxref_22_1 N_MM3_g 0.00183957f
cc_141 N_noxref_22_1 N_CLKB_6 0.000104327f
cc_142 N_noxref_22_1 N_CLKB_18 0.000551242f
cc_143 N_noxref_22_1 N_noxref_20_1 0.0076875f
cc_144 N_noxref_22_1 N_noxref_21_1 0.000463746f
x_PM_DFFHQNx3_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_DFFHQNx3_ASAP7_75t_R%noxref_23
cc_145 N_noxref_23_1 N_MM3_g 0.00185344f
cc_146 N_noxref_23_1 N_CLKB_7 0.000100593f
cc_147 N_noxref_23_1 N_CLKB_19 0.000556726f
cc_148 N_noxref_23_1 N_noxref_20_1 0.000463573f
cc_149 N_noxref_23_1 N_noxref_21_1 0.00769135f
cc_150 N_noxref_23_1 N_noxref_22_1 0.00122173f
x_PM_DFFHQNx3_ASAP7_75t_R%PD2 VSS N_MM10_s N_MM11_d N_PD2_4 N_PD2_5 N_PD2_1
+ PM_DFFHQNx3_ASAP7_75t_R%PD2
cc_151 N_PD2_4 N_MM10_g 0.0150485f
cc_152 N_PD2_5 N_CLKB_8 0.0014696f
cc_153 N_PD2_1 N_CLKB_2 0.000539911f
cc_154 N_PD2_1 N_MM9_g 0.00206219f
cc_155 N_PD2_4 N_MM9_g 0.00714091f
cc_156 N_PD2_5 N_MM9_g 0.024057f
cc_157 N_PD2_5 N_MM11_g 0.0146029f
cc_158 N_PD2_1 N_MH_14 0.000435677f
cc_159 N_PD2_4 N_MH_3 0.00061455f
cc_160 N_PD2_1 N_MH_20 0.00320686f
x_PM_DFFHQNx3_ASAP7_75t_R%SS VSS N_MM19_g N_MM14_d N_MM15_d N_SS_12 N_SS_10
+ N_SS_11 N_SS_15 N_SS_4 N_SS_3 N_SS_14 N_SS_1 N_SS_16 N_SS_13
+ PM_DFFHQNx3_ASAP7_75t_R%SS
cc_161 N_MM19_g N_CLKB_8 0.000215376f
cc_162 N_MM19_g N_CLKB_4 0.000537906f
cc_163 N_MM19_g N_MM18_g 0.0135403f
x_PM_DFFHQNx3_ASAP7_75t_R%MS VSS N_MM11_g N_MM6_d N_MM12_d N_MM7_d N_MM13_d
+ N_MS_13 N_MS_17 N_MS_18 N_MS_14 N_MS_3 N_MS_15 N_MS_12 N_MS_1 N_MS_11 N_MS_4
+ N_MS_16 PM_DFFHQNx3_ASAP7_75t_R%MS
cc_164 N_MS_13 N_MM10_g 0.000130138f
cc_165 N_MS_13 N_CLKN_24 0.000324163f
cc_166 N_MS_13 N_CLKN_28 0.00022929f
cc_167 N_MS_13 N_CLKN_3 0.000229581f
cc_168 N_MS_17 N_CLKN_24 0.00452644f
cc_169 N_MS_17 N_CLKN_3 0.000282384f
cc_170 N_MS_18 N_CLKN_24 0.000632715f
cc_171 N_MS_14 N_CLKN_28 0.0027899f
cc_172 N_MS_13 N_MM13_g 0.0153408f
cc_173 N_MS_3 N_CLKB_8 0.00055579f
cc_174 N_MS_3 N_CLKB_2 0.000123737f
cc_175 N_MS_3 N_CLKB_22 0.000157903f
cc_176 N_MS_3 N_MM9_g 0.000165533f
cc_177 N_MS_3 N_CLKB_26 0.000172147f
cc_178 N_MS_15 N_CLKB_22 0.000290783f
cc_179 N_MS_12 N_MM12_g 0.0078041f
cc_180 N_MS_13 N_MM12_g 0.00777346f
cc_181 N_MS_15 N_CLKB_8 0.000383383f
cc_182 N_MS_1 N_MM9_g 0.000560232f
cc_183 N_MS_17 N_CLKB_8 0.00157508f
cc_184 N_MS_11 N_MM12_g 0.00651789f
cc_185 N_MS_4 N_MM12_g 0.00255242f
cc_186 N_MS_4 N_CLKB_8 0.00635858f
cc_187 N_MM11_g N_MM9_g 0.0142057f
cc_188 N_MS_3 N_MM12_g 0.0259348f
x_PM_DFFHQNx3_ASAP7_75t_R%CLKB VSS N_MM1_g N_MM9_g N_MM12_g N_MM18_g N_MM23_d
+ N_MM22_d N_CLKB_18 N_CLKB_20 N_CLKB_26 N_CLKB_6 N_CLKB_7 N_CLKB_23 N_CLKB_24
+ N_CLKB_4 N_CLKB_25 N_CLKB_22 N_CLKB_19 N_CLKB_1 N_CLKB_21 N_CLKB_8 N_CLKB_2
+ PM_DFFHQNx3_ASAP7_75t_R%CLKB
cc_189 N_CLKB_18 N_CLK_6 8.57854e-20
cc_190 N_CLKB_20 N_CLK_6 9.12674e-20
cc_191 N_CLKB_26 N_CLK_6 0.000123342f
cc_192 N_CLKB_6 N_CLK_6 0.000361693f
cc_193 N_CLKB_7 N_CLK_6 0.000387298f
cc_194 N_CLKB_23 N_CLK_7 0.000500038f
cc_195 N_CLKB_20 N_CLK_8 0.000514675f
cc_196 N_CLKB_23 N_CLK_5 0.00120151f
cc_197 N_CLKB_24 N_CLK_6 0.00199622f
cc_198 N_CLKB_6 N_MM22_g 0.000721222f
cc_199 N_CLKB_7 N_MM22_g 0.000747071f
cc_200 N_CLKB_4 N_MM13_g 0.000222558f
cc_201 N_CLKB_25 N_CLKN_28 0.000285919f
cc_202 N_CLKB_22 N_CLKN_28 0.000669652f
cc_203 N_CLKB_24 N_CLKN_22 0.000310766f
cc_204 N_CLKB_19 N_MM22_g 0.0110945f
cc_205 N_CLKB_23 N_CLKN_22 0.000357496f
cc_206 N_CLKB_1 N_CLKN_2 0.00169517f
cc_207 N_CLKB_21 N_CLKN_28 0.00104596f
cc_208 N_CLKB_20 N_CLKN_22 0.00766547f
cc_209 N_CLKB_20 N_CLKN_28 0.000519084f
cc_210 N_CLKB_8 N_CLKN_24 0.000534461f
cc_211 N_CLKB_25 N_CLKN_2 0.000549016f
cc_212 N_CLKB_2 N_MM10_g 0.000589093f
cc_213 N_CLKB_26 N_CLKN_23 0.000616959f
cc_214 N_CLKB_8 N_CLKN_3 0.00279616f
cc_215 N_CLKB_20 N_CLKN_1 0.000691464f
cc_216 N_CLKB_19 N_CLKN_1 0.00121517f
cc_217 N_MM1_g N_MM10_g 0.00163577f
cc_218 N_CLKB_25 N_CLKN_23 0.00263609f
cc_219 N_CLKB_8 N_MM13_g 0.00423843f
cc_220 N_MM12_g N_MM13_g 0.00572282f
cc_221 N_MM9_g N_MM10_g 0.00910623f
cc_222 N_MM18_g N_MM13_g 0.0184454f
cc_223 N_CLKB_26 N_CLKN_28 0.031089f
cc_224 N_CLKB_18 N_MM22_g 0.038903f
cc_225 N_CLKB_6 N_MM3_g 0.00011685f
cc_226 N_CLKB_21 N_MM3_g 0.000132909f
cc_227 N_CLKB_20 N_MM3_g 0.000186961f
cc_228 N_CLKB_1 N_MM3_g 0.000265584f
cc_229 N_CLKB_25 N_MM3_g 0.000617636f
cc_230 N_CLKB_23 N_D_7 0.000843543f
cc_231 N_CLKB_26 N_D_6 0.00108916f
cc_232 N_CLKB_21 N_D_6 0.0011142f
cc_233 N_CLKB_24 N_D_9 0.00121817f
cc_234 N_CLKB_1 N_D_1 0.00161854f
cc_235 N_CLKB_20 N_D_4 0.00180998f
cc_236 N_CLKB_25 N_D_6 0.00203563f
cc_237 N_CLKB_20 N_D_5 0.00266241f
cc_238 N_CLKB_20 N_D_8 0.00411749f
cc_239 N_MM1_g N_MM3_g 0.00527306f
x_PM_DFFHQNx3_ASAP7_75t_R%SH VSS N_MM14_g N_MM24_g N_MM24@3_g N_MM24@2_g
+ N_MM13_s N_MM18_d N_MM12_s N_MM17_d N_SH_30 N_SH_6 N_SH_20 N_SH_16 N_SH_15
+ N_SH_25 N_SH_27 N_SH_18 N_SH_19 N_SH_17 N_SH_5 N_SH_23 N_SH_29 N_SH_2 N_SH_28
+ N_SH_24 N_SH_22 N_SH_1 N_SH_26 N_SH_21 PM_DFFHQNx3_ASAP7_75t_R%SH
cc_240 N_SH_30 N_CLKN_28 0.000137532f
cc_241 N_SH_6 N_MM13_g 0.000163831f
cc_242 N_SH_20 N_CLKN_24 0.000212662f
cc_243 N_SH_16 N_MM13_g 0.00675259f
cc_244 N_SH_15 N_MM13_g 0.0067885f
cc_245 N_SH_25 N_CLKN_24 0.000353729f
cc_246 N_SH_27 N_CLKN_24 0.000935658f
cc_247 N_SH_18 N_CLKN_3 0.000445115f
cc_248 N_SH_19 N_CLKN_24 0.000522982f
cc_249 N_SH_17 N_CLKN_24 0.000529757f
cc_250 N_SH_5 N_CLKN_3 0.000536728f
cc_251 N_SH_17 N_CLKN_28 0.00111054f
cc_252 N_SH_18 N_CLKN_24 0.00388722f
cc_253 N_SH_5 N_MM13_g 0.0184293f
cc_254 N_SH_17 N_CLKB_26 9.11347e-20
cc_255 N_SH_25 N_CLKB_8 0.000184575f
cc_256 N_SH_27 N_CLKB_8 0.000201135f
cc_257 N_SH_15 N_MM12_g 0.00677653f
cc_258 N_SH_6 N_CLKB_8 0.000297547f
cc_259 N_SH_20 N_CLKB_4 0.000403199f
cc_260 N_SH_18 N_CLKB_8 0.000420117f
cc_261 N_SH_19 N_CLKB_8 0.000613345f
cc_262 N_SH_16 N_CLKB_4 0.000928311f
cc_263 N_SH_6 N_MM18_g 0.000989101f
cc_264 N_SH_16 N_CLKB_8 0.00230339f
cc_265 N_SH_5 N_MM12_g 0.00951501f
cc_266 N_SH_16 N_MM18_g 0.016274f
cc_267 N_SH_19 N_MS_3 9.71132e-20
cc_268 N_SH_18 N_MS_3 0.000112268f
cc_269 N_SH_25 N_MS_3 0.00013281f
cc_270 N_SH_6 N_MS_3 0.000211236f
cc_271 N_SH_16 N_MS_3 0.000438565f
cc_272 N_SH_15 N_MS_3 0.000463915f
cc_273 N_SH_25 N_MS_4 0.000318288f
cc_274 N_SH_6 N_MS_4 0.000418085f
cc_275 N_SH_17 N_MS_16 0.000525587f
cc_276 N_SH_16 N_MS_4 0.000582695f
cc_277 N_SH_25 N_MS_17 0.000616175f
cc_278 N_SH_17 N_MS_18 0.00165552f
cc_279 N_SH_5 N_MS_3 0.00369603f
cc_280 N_SH_17 N_MM19_g 9.54229e-20
cc_281 N_SH_23 N_MM19_g 0.000129092f
cc_282 N_SH_19 N_MM19_g 0.000140302f
cc_283 N_SH_29 N_MM19_g 0.00018262f
cc_284 N_SH_2 N_MM19_g 0.000194841f
cc_285 N_SH_28 N_SS_12 0.000215496f
cc_286 N_MM14_g N_SS_10 0.00686379f
cc_287 N_MM14_g N_SS_11 0.00682988f
cc_288 N_SH_2 N_SS_15 0.000280575f
cc_289 N_SH_24 N_SS_15 0.00631225f
cc_290 N_SH_22 N_SS_4 0.000330589f
cc_291 N_MM14_g N_SS_3 0.000397637f
cc_292 N_SH_23 N_SS_15 0.00186396f
cc_293 N_MM14_g N_SS_4 0.000516529f
cc_294 N_SH_22 N_SS_14 0.000651121f
cc_295 N_SH_1 N_SS_1 0.000686419f
cc_296 N_SH_26 N_SS_16 0.000794357f
cc_297 N_SH_18 N_SS_1 0.000849146f
cc_298 N_SH_29 N_SS_15 0.000900846f
cc_299 N_SH_21 N_SS_12 0.000945454f
cc_300 N_SH_23 N_SS_13 0.0010905f
cc_301 N_MM14_g N_SS_1 0.00113556f
cc_302 N_SH_29 N_SS_14 0.00128145f
cc_303 N_SH_1 N_MM19_g 0.00129777f
cc_304 N_SH_20 N_SS_12 0.00152066f
cc_305 N_SH_30 N_SS_15 0.00187742f
cc_306 N_SH_18 N_SS_12 0.00470692f
cc_307 N_MM14_g N_MM19_g 0.0293467f
x_PM_DFFHQNx3_ASAP7_75t_R%CLKN VSS N_MM22_g N_MM10_g N_MM13_g N_MM20_d N_MM21_d
+ N_CLKN_22 N_CLKN_8 N_CLKN_26 N_CLKN_7 N_CLKN_16 N_CLKN_17 N_CLKN_1 N_CLKN_19
+ N_CLKN_21 N_CLKN_20 N_CLKN_18 N_CLKN_28 N_CLKN_23 N_CLKN_2 N_CLKN_24 N_CLKN_3
+ PM_DFFHQNx3_ASAP7_75t_R%CLKN
cc_308 N_CLKN_22 N_MM20_g 0.000243475f
cc_309 N_CLKN_8 N_MM20_g 0.00112888f
cc_310 N_CLKN_26 N_MM20_g 0.000252097f
cc_311 N_CLKN_7 N_MM20_g 0.0011647f
cc_312 N_CLKN_16 N_MM20_g 0.0112193f
cc_313 N_CLKN_17 N_MM20_g 0.0113277f
cc_314 N_CLKN_1 N_CLK_8 0.000441582f
cc_315 N_CLKN_19 N_CLK_8 0.000504575f
cc_316 N_CLKN_21 N_CLK_8 0.000765329f
cc_317 N_CLKN_20 N_CLK_5 0.000800078f
cc_318 N_CLKN_26 N_CLK_1 0.000803931f
cc_319 N_CLKN_21 N_CLK_6 0.000842599f
cc_320 N_CLKN_22 N_CLK_7 0.001063f
cc_321 N_CLKN_18 N_CLK_7 0.00116394f
cc_322 N_CLKN_28 N_CLK_8 0.00178169f
cc_323 N_CLKN_26 N_CLK_8 0.00178252f
cc_324 N_CLKN_1 N_CLK_1 0.00248534f
cc_325 N_CLKN_20 N_CLK_7 0.00268142f
cc_326 N_CLKN_22 N_CLK_8 0.00324624f
cc_327 N_CLKN_26 N_CLK_4 0.00343261f
cc_328 N_MM22_g N_MM20_g 0.0350536f
*END of DFFHQNx3_ASAP7_75t_R.pxi
.ENDS
** Design:	DFFHQx4_ASAP7_75t_R
* Created:	"Fri Aug 17 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "DFFHQx4_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "DFFHQx4_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_DFFHQx4_ASAP7_75t_R%noxref_29 VSS 1
c1 1 VSS 0.0422386f
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%noxref_30 VSS 1
c1 1 VSS 0.0422877f
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%Q VSS 35 26 27 41 42 50 51 54 55 14 18 16 15 13
+ 21 20 2 3 4 1
c1 1 VSS 0.00896302f
c2 2 VSS 0.00876961f
c3 3 VSS 0.00949415f
c4 4 VSS 0.010041f
c5 13 VSS 0.00449514f
c6 14 VSS 0.00445213f
c7 15 VSS 0.00444851f
c8 16 VSS 0.00439519f
c9 17 VSS 0.0167002f
c10 18 VSS 0.0170325f
c11 19 VSS 0.00775503f
c12 20 VSS 0.00288792f
c13 21 VSS 0.00342737f
c14 22 VSS 0.00326848f
c15 23 VSS 0.00324858f
r1 55 53 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.1510 $Y=0.2025 $X2=1.1485 $Y2=0.2025
r2 2 53 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.1340 $Y=0.2025 $X2=1.1485 $Y2=0.2025
r3 15 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.1195 $Y=0.2025 $X2=1.1340 $Y2=0.2025
r4 54 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.1170 $Y=0.2025 $X2=1.1195 $Y2=0.2025
r5 2 47 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.1340 $Y=0.2025
+ $X2=1.1340 $Y2=0.2160
r6 51 49 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.2590 $Y=0.2025 $X2=1.2565 $Y2=0.2025
r7 4 49 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.2420 $Y=0.2025 $X2=1.2565 $Y2=0.2025
r8 16 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.2275 $Y=0.2025 $X2=1.2420 $Y2=0.2025
r9 50 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.2250 $Y=0.2025 $X2=1.2275 $Y2=0.2025
r10 21 45 4.64944 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.1340
+ $Y=0.2340 $X2=1.1590 $Y2=0.2340
r11 21 47 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.1340
+ $Y=0.2340 $X2=1.1340 $Y2=0.2160
r12 4 43 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.2420 $Y=0.2025
+ $X2=1.2420 $Y2=0.2340
r13 43 44 9.32759 $w=1.3e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=1.2420
+ $Y=0.2340 $X2=1.2820 $Y2=0.2340
r14 18 43 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.2040
+ $Y=0.2340 $X2=1.2420 $Y2=0.2340
r15 18 45 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.2040
+ $Y=0.2340 $X2=1.1590 $Y2=0.2340
r16 23 38 2.48126 $w=1.71429e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3230 $Y=0.2340 $X2=1.3230 $Y2=0.2130
r17 23 44 7.66726 $w=1.56829e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3230 $Y=0.2340 $X2=1.2820 $Y2=0.2340
r18 42 40 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.2590 $Y=0.0675 $X2=1.2565 $Y2=0.0675
r19 3 40 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.2420 $Y=0.0675 $X2=1.2565 $Y2=0.0675
r20 14 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.2275 $Y=0.0675 $X2=1.2420 $Y2=0.0675
r21 41 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.2250 $Y=0.0675 $X2=1.2275 $Y2=0.0675
r22 37 38 6.8096 $w=1.5e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.1730 $X2=1.3230 $Y2=0.2130
r23 36 37 5.66048 $w=1.5e-08 $l=3.33e-08 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.1397 $X2=1.3230 $Y2=0.1730
r24 35 36 0.97888 $w=1.5e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.1340 $X2=1.3230 $Y2=0.1397
r25 35 34 0.6384 $w=1.5e-08 $l=3.8e-09 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.1340 $X2=1.3230 $Y2=0.1302
r26 33 34 5.49024 $w=1.5e-08 $l=3.22e-08 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.0980 $X2=1.3230 $Y2=0.1302
r27 19 22 2.48126 $w=1.71429e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3230 $Y=0.0570 $X2=1.3230 $Y2=0.0360
r28 19 33 6.97984 $w=1.5e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.0570 $X2=1.3230 $Y2=0.0980
r29 3 31 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.2420 $Y=0.0675
+ $X2=1.2420 $Y2=0.0360
r30 22 32 7.66726 $w=1.56829e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3230 $Y=0.0360 $X2=1.2820 $Y2=0.0360
r31 31 32 9.32759 $w=1.3e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=1.2420
+ $Y=0.0360 $X2=1.2820 $Y2=0.0360
r32 30 31 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.2040
+ $Y=0.0360 $X2=1.2420 $Y2=0.0360
r33 17 29 4.64944 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.1590
+ $Y=0.0360 $X2=1.1340 $Y2=0.0360
r34 17 30 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.1590
+ $Y=0.0360 $X2=1.2040 $Y2=0.0360
r35 20 29 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.1340
+ $Y=0.0540 $X2=1.1340 $Y2=0.0360
r36 1 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.1340 $Y=0.0675
+ $X2=1.1340 $Y2=0.0540
r37 27 25 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.1510 $Y=0.0675 $X2=1.1485 $Y2=0.0675
r38 1 25 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.1340 $Y=0.0675 $X2=1.1485 $Y2=0.0675
r39 13 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.1195 $Y=0.0675 $X2=1.1340 $Y2=0.0675
r40 26 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.1170 $Y=0.0675 $X2=1.1195 $Y2=0.0675
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%PD3 VSS 2 4 1
c1 1 VSS 0.00097274f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0405 $X2=0.4905 $Y2=0.0405
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0405 $X2=0.4735 $Y2=0.0405
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4735 $Y=0.0405 $X2=0.4905 $Y2=0.0405
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.0415651f
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%PD4 VSS 2 4 1
c1 1 VSS 0.000952912f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.2295 $X2=0.7605 $Y2=0.2295
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.2295 $X2=0.7435 $Y2=0.2295
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7435 $Y=0.2295 $X2=0.7605 $Y2=0.2295
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%PU1 VSS 2 4 1
c1 1 VSS 0.000988923f
r1 4 3 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3365 $Y2=0.2025
r2 2 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3195 $Y2=0.2025
r3 1 3 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3195 $Y=0.2025 $X2=0.3365 $Y2=0.2025
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.0415489f
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.00491256f
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.004928f
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%D VSS 19 3 5 6 7 9 1 4 8
c1 1 VSS 0.0109493f
c2 3 VSS 0.0835668f
c3 4 VSS 0.003706f
c4 5 VSS 0.00336744f
c5 6 VSS 0.00165307f
c6 7 VSS 0.00749114f
c7 8 VSS 0.00108235f
c8 9 VSS 0.00643786f
r1 9 21 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2430 $Y2=0.2140
r2 7 18 5.17411 $w=1.46514e-08 $l=2.72e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0360 $X2=0.2430 $Y2=0.0632
r3 5 8 7.7975 $w=1.41688e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1735 $X2=0.2430 $Y2=0.1350
r4 5 21 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1735 $X2=0.2430 $Y2=0.2140
r5 19 20 2.85657 $w=1.3e-08 $l=1.22e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0820 $X2=0.2430 $Y2=0.0942
r6 19 18 4.37231 $w=1.3e-08 $l=1.88e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0820 $X2=0.2430 $Y2=0.0632
r7 4 8 3.2503 $w=1.53684e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1160 $X2=0.2430 $Y2=0.1350
r8 4 20 5.07188 $w=1.3e-08 $l=2.18e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1160 $X2=0.2430 $Y2=0.0942
r9 16 17 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2715
+ $Y=0.1350 $X2=0.2810 $Y2=0.1350
r10 6 16 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2615
+ $Y=0.1350 $X2=0.2715 $Y2=0.1350
r11 6 8 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2615 $Y=0.1350 $X2=0.2430 $Y2=0.1350
r12 14 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2770 $Y=0.1350
+ $X2=0.2810 $Y2=0.1350
r13 12 14 4.43042 $w=1.53e-08 $l=7.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.2845 $Y=0.1350 $X2=0.2770 $Y2=0.1350
r14 1 11 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.2885
+ $Y=0.1350 $X2=0.2985 $Y2=0.1350
r15 1 12 1.86855 $w=1.78125e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.2885 $Y=0.1350 $X2=0.2845 $Y2=0.1350
r16 3 11 2.53453 $w=1.32811e-07 $l=1.5e-09 $layer=LIG $thickness=5.23243e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2985 $Y2=0.1350
r17 3 12 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2845 $Y2=0.1350
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%noxref_26 VSS 1
c1 1 VSS 0.00423748f
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%noxref_28 VSS 1
c1 1 VSS 0.0415404f
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%noxref_27 VSS 1
c1 1 VSS 0.0415022f
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.00421725f
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%SS VSS 9 31 41 10 11 4 15 3 14 1 16 12 13
c1 1 VSS 0.00117155f
c2 3 VSS 0.00611629f
c3 4 VSS 0.00666211f
c4 9 VSS 0.0384353f
c5 10 VSS 0.00320705f
c6 11 VSS 0.00319459f
c7 12 VSS 0.0019451f
c8 13 VSS 0.013056f
c9 14 VSS 0.00918443f
c10 15 VSS 0.00755396f
c11 16 VSS 0.00269165f
c12 17 VSS 0.00421963f
c13 18 VSS 0.00366179f
r1 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.2295 $X2=0.8620 $Y2=0.2295
r2 41 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.2295 $X2=0.8495 $Y2=0.2295
r3 4 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.2295
+ $X2=0.8640 $Y2=0.2340
r4 38 39 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.2340 $X2=0.8865 $Y2=0.2340
r5 14 18 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9180 $Y=0.2340 $X2=0.9450 $Y2=0.2340
r6 14 39 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.2340 $X2=0.8865 $Y2=0.2340
r7 18 36 0.56619 $w=2.22842e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.2340 $X2=0.9450 $Y2=0.2245
r8 35 36 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1975 $X2=0.9450 $Y2=0.2245
r9 34 35 6.64591 $w=1.3e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1690 $X2=0.9450 $Y2=0.1975
r10 33 34 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1445 $X2=0.9450 $Y2=0.1690
r11 32 33 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1195 $X2=0.9450 $Y2=0.1445
r12 15 17 8.84443 $w=1.496e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.0810 $X2=0.9450 $Y2=0.0360
r13 15 32 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.0810 $X2=0.9450 $Y2=0.1195
r14 10 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.0405 $X2=0.8620 $Y2=0.0405
r15 31 10 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.0405 $X2=0.8495 $Y2=0.0405
r16 17 29 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.0360 $X2=0.9180 $Y2=0.0360
r17 3 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.0405
+ $X2=0.8640 $Y2=0.0360
r18 28 29 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.0360 $X2=0.9180 $Y2=0.0360
r19 27 28 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.0360 $X2=0.8910 $Y2=0.0360
r20 26 27 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.0360 $X2=0.8640 $Y2=0.0360
r21 13 16 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.0360 $X2=0.7830 $Y2=0.0360
r22 13 26 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0360 $X2=0.8370 $Y2=0.0360
r23 12 23 8.04505 $w=1.3e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.0705 $X2=0.7830 $Y2=0.1050
r24 12 16 6.39593 $w=1.55565e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7830 $Y=0.0705 $X2=0.7830 $Y2=0.0360
r25 1 20 2.36633 $w=2.3e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.7830
+ $Y=0.1055 $X2=0.7830 $Y2=0.1055
r26 1 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7830 $Y=0.1055
+ $X2=0.7830 $Y2=0.1050
r27 9 20 0.314665 $w=2.27e-07 $l=2.95e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.7830 $Y=0.1350 $X2=0.7830 $Y2=0.1055
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%PD5 VSS 7 12 4 1 5
c1 1 VSS 0.00736396f
c2 4 VSS 0.00187625f
c3 5 VSS 0.00237272f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.0405 $X2=0.7705 $Y2=0.0405
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7580 $Y=0.0405 $X2=0.7705 $Y2=0.0405
r3 9 5 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.7425
+ $Y=0.0405 $X2=0.7560 $Y2=0.0405
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.7275
+ $Y=0.0405 $X2=0.7425 $Y2=0.0405
r5 1 8 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.7020
+ $Y=0.0405 $X2=0.7275 $Y2=0.0405
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.0405 $X2=0.7000 $Y2=0.0405
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.0405 $X2=0.6875 $Y2=0.0405
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%NET049 VSS 9 10 11 12 62 63 66 67 13 16 4 17 18
+ 14 3 1 22 20 19
c1 1 VSS 0.0190246f
c2 3 VSS 0.0132034f
c3 4 VSS 0.0137464f
c4 9 VSS 0.0817164f
c5 10 VSS 0.0814408f
c6 11 VSS 0.0816409f
c7 12 VSS 0.0820926f
c8 13 VSS 0.00823027f
c9 14 VSS 0.00822518f
c10 15 VSS 0.00924619f
c11 16 VSS 0.00861171f
c12 17 VSS 0.00393415f
c13 18 VSS 0.00383151f
c14 19 VSS 0.00289129f
c15 20 VSS 0.00432644f
c16 21 VSS 0.00142877f
c17 22 VSS 0.00355378f
r1 67 65 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0430 $Y=0.2025 $X2=1.0405 $Y2=0.2025
r2 4 65 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0260 $Y=0.2025 $X2=1.0405 $Y2=0.2025
r3 14 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0115 $Y=0.2025 $X2=1.0260 $Y2=0.2025
r4 66 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0090 $Y=0.2025 $X2=1.0115 $Y2=0.2025
r5 63 61 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.0430 $Y=0.0675 $X2=1.0405 $Y2=0.0675
r6 3 61 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.0260 $Y=0.0675 $X2=1.0405 $Y2=0.0675
r7 13 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.0115 $Y=0.0675 $X2=1.0260 $Y2=0.0675
r8 62 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.0090 $Y=0.0675 $X2=1.0115 $Y2=0.0675
r9 4 58 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0260 $Y=0.2025
+ $X2=1.0260 $Y2=0.2340
r10 3 56 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0260 $Y=0.0675
+ $X2=1.0260 $Y2=0.0360
r11 58 59 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.2340 $X2=1.0575 $Y2=0.2340
r12 16 58 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.0145
+ $Y=0.2340 $X2=1.0260 $Y2=0.2340
r13 56 57 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.0360 $X2=1.0575 $Y2=0.0360
r14 15 56 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.0145
+ $Y=0.0360 $X2=1.0260 $Y2=0.0360
r15 22 55 3.24787 $w=1.72e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.0890
+ $Y=0.2340 $X2=1.0890 $Y2=0.2130
r16 22 59 5.69637 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0890 $Y=0.2340 $X2=1.0575 $Y2=0.2340
r17 20 53 3.24787 $w=1.72e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.0890
+ $Y=0.0360 $X2=1.0890 $Y2=0.0570
r18 20 57 5.69637 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0890 $Y=0.0360 $X2=1.0575 $Y2=0.0360
r19 54 55 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=1.0890
+ $Y=0.1840 $X2=1.0890 $Y2=0.2130
r20 18 21 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=1.0890
+ $Y=0.1560 $X2=1.0890 $Y2=0.1360
r21 18 54 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.0890
+ $Y=0.1560 $X2=1.0890 $Y2=0.1840
r22 52 53 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=1.0890
+ $Y=0.0955 $X2=1.0890 $Y2=0.0570
r23 17 21 1.50137 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0890 $Y=0.1245 $X2=1.0890 $Y2=0.1360
r24 17 52 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=1.0890
+ $Y=0.1245 $X2=1.0890 $Y2=0.0955
r25 21 49 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.0890
+ $Y=0.1360 $X2=1.1115 $Y2=0.1360
r26 12 43 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=1.2690
+ $Y=0.1350 $X2=1.2690 $Y2=0.1360
r27 11 37 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=1.2150
+ $Y=0.1350 $X2=1.2150 $Y2=0.1360
r28 48 49 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.1340
+ $Y=0.1360 $X2=1.1115 $Y2=0.1360
r29 19 46 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.1475
+ $Y=0.1360 $X2=1.1610 $Y2=0.1360
r30 19 48 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.1475
+ $Y=0.1360 $X2=1.1340 $Y2=0.1360
r31 10 30 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=1.1610 $Y=0.1350 $X2=1.1610 $Y2=0.1360
r32 41 43 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.2565 $Y=0.1360 $X2=1.2690 $Y2=0.1360
r33 40 41 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.2420 $Y=0.1360 $X2=1.2565 $Y2=0.1360
r34 38 40 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.2275 $Y=0.1360 $X2=1.2420 $Y2=0.1360
r35 37 38 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.2150 $Y=0.1360 $X2=1.2275 $Y2=0.1360
r36 35 37 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.2025 $Y=0.1360 $X2=1.2150 $Y2=0.1360
r37 34 35 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.1880 $Y=0.1360 $X2=1.2025 $Y2=0.1360
r38 32 34 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.1735 $Y=0.1360 $X2=1.1880 $Y2=0.1360
r39 31 32 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=1.1705 $Y=0.1360 $X2=1.1735 $Y2=0.1360
r40 30 31 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=1.1610
+ $Y=0.1360 $X2=1.1705 $Y2=0.1360
r41 30 46 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.1610 $Y=0.1360
+ $X2=1.1610 $Y2=0.1360
r42 29 30 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=1.1515
+ $Y=0.1360 $X2=1.1610 $Y2=0.1360
r43 27 29 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=1.1485 $Y=0.1360 $X2=1.1515 $Y2=0.1360
r44 26 27 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.1340 $Y=0.1360 $X2=1.1485 $Y2=0.1360
r45 25 26 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.1195 $Y=0.1360 $X2=1.1340 $Y2=0.1360
r46 9 1 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=1.1070
+ $Y=0.1350 $X2=1.1070 $Y2=0.1360
r47 1 24 2.90696 $w=2.1681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.1070 $Y=0.1360 $X2=1.0965 $Y2=0.1360
r48 1 25 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.1070 $Y=0.1360 $X2=1.1195 $Y2=0.1360
r49 9 24 0.610027 $w=2.16919e-07 $l=1.05475e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=1.1070 $Y=0.1350 $X2=1.0965 $Y2=0.1360
r50 9 25 1.79147 $w=1.8466e-07 $l=1.25399e-08 $layer=LIG $thickness=5.44e-08
+ $X=1.1070 $Y=0.1350 $X2=1.1195 $Y2=0.1360
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%SH VSS 11 12 13 74 77 81 84 5 6 19 14 15 24 26
+ 17 18 16 22 2 28 27 21 23 1 25 20 29
c1 1 VSS 0.000781112f
c2 2 VSS 0.00780299f
c3 5 VSS 0.00511021f
c4 6 VSS 0.00487233f
c5 11 VSS 0.0374674f
c6 12 VSS 0.081032f
c7 13 VSS 0.0809455f
c8 14 VSS 0.00498732f
c9 15 VSS 0.00519827f
c10 16 VSS 0.00840732f
c11 17 VSS 0.00193507f
c12 18 VSS 0.0018376f
c13 19 VSS 0.00259979f
c14 20 VSS 0.000803918f
c15 21 VSS 0.000473119f
c16 22 VSS 0.0013086f
c17 23 VSS 0.00262965f
c18 24 VSS 0.00659022f
c19 25 VSS 0.00266206f
c20 26 VSS 0.000112382f
c21 27 VSS 0.000394971f
c22 28 VSS 0.000377583f
c23 29 VSS 0.00987851f
r1 84 83 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r2 5 83 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6500 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r3 80 5 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6380 $Y=0.0405 $X2=0.6500 $Y2=0.0405
r4 14 80 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0405 $X2=0.6380 $Y2=0.0405
r5 81 14 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.0405 $X2=0.6335 $Y2=0.0405
r6 13 68 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=1.0530
+ $Y=0.1350 $X2=1.0530 $Y2=0.1360
r7 12 60 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.9990 $Y=0.1350 $X2=0.9990 $Y2=0.1360
r8 77 76 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r9 75 76 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7120 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r10 6 75 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7000 $Y=0.2295 $X2=0.7120 $Y2=0.2295
r11 15 6 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.2295 $X2=0.7000 $Y2=0.2295
r12 74 15 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.2295 $X2=0.6875 $Y2=0.2295
r13 5 58 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.0405
+ $X2=0.6480 $Y2=0.0360
r14 66 68 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.0405 $Y=0.1360 $X2=1.0530 $Y2=0.1360
r15 65 66 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.0260 $Y=0.1360 $X2=1.0405 $Y2=0.1360
r16 63 65 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.0115 $Y=0.1360 $X2=1.0260 $Y2=0.1360
r17 61 63 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=1.0085 $Y=0.1360 $X2=1.0115 $Y2=0.1360
r18 60 61 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.9990
+ $Y=0.1360 $X2=1.0085 $Y2=0.1360
r19 2 60 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.9895
+ $Y=0.1360 $X2=0.9990 $Y2=0.1360
r20 6 51 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7020 $Y=0.2295
+ $X2=0.7020 $Y2=0.2330
r21 58 59 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6480
+ $Y=0.0360 $X2=0.6615 $Y2=0.0360
r22 56 59 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0360 $X2=0.6615 $Y2=0.0360
r23 55 56 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6860
+ $Y=0.0360 $X2=0.6750 $Y2=0.0360
r24 16 25 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.7040
+ $Y=0.0360 $X2=0.7290 $Y2=0.0360
r25 16 55 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7040
+ $Y=0.0360 $X2=0.6860 $Y2=0.0360
r26 53 60 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.9990 $Y=0.1445
+ $X2=0.9990 $Y2=0.1360
r27 23 53 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.9990
+ $Y=0.1245 $X2=0.9990 $Y2=0.1445
r28 51 52 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.2330 $X2=0.7155 $Y2=0.2330
r29 24 52 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.2330 $X2=0.7155 $Y2=0.2330
r30 25 44 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.0360 $X2=0.7290 $Y2=0.0630
r31 48 53 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.9990 $Y=0.1530
+ $X2=0.9990 $Y2=0.1445
r32 47 48 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1530 $X2=0.9990 $Y2=0.1530
r33 46 47 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1530 $X2=0.9450 $Y2=0.1530
r34 29 46 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.8795
+ $Y=0.1530 $X2=0.8910 $Y2=0.1530
r35 45 46 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.8910 $Y=0.1485 $X2=0.8910
+ $Y2=0.1530
r36 22 45 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1305 $X2=0.8910 $Y2=0.1485
r37 18 39 6.38362 $w=1.33509e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1975 $X2=0.7290 $Y2=0.1690
r38 18 24 7.09793 $w=1.42676e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1975 $X2=0.7290 $Y2=0.2330
r39 43 44 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.0900 $X2=0.7290 $Y2=0.0630
r40 42 43 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1000 $X2=0.7290 $Y2=0.0900
r41 41 42 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1100 $X2=0.7290 $Y2=0.1000
r42 17 26 4.67854 $w=1.44583e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1360 $X2=0.7290 $Y2=0.1600
r43 17 41 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1360 $X2=0.7290 $Y2=0.1100
r44 28 40 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1575 $X2=0.8910 $Y2=0.1665
r45 28 45 1.50855 $w=1.55e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1575 $X2=0.8910 $Y2=0.1485
r46 28 46 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.8910 $Y=0.1575 $X2=0.8910
+ $Y2=0.1530
r47 26 39 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1600 $X2=0.7290 $Y2=0.1690
r48 38 40 4.19024 $w=1.156e-08 $l=2.54018e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8660 $Y=0.1620 $X2=0.8910 $Y2=0.1665
r49 21 27 1.38478 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8480 $Y=0.1620 $X2=0.8370 $Y2=0.1620
r50 21 38 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8480
+ $Y=0.1620 $X2=0.8660 $Y2=0.1620
r51 37 39 4.4015 $w=1.35e-08 $l=2.78927e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7560 $Y=0.1620 $X2=0.7290 $Y2=0.1690
r52 36 37 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1620 $X2=0.7560 $Y2=0.1620
r53 19 27 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.1620 $X2=0.8370 $Y2=0.1620
r54 19 36 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.1620 $X2=0.7830 $Y2=0.1620
r55 27 35 4.88263 $w=1.47308e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8370 $Y=0.1620 $X2=0.8370 $Y2=0.1360
r56 20 35 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1180 $X2=0.8370 $Y2=0.1360
r57 11 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.8370
+ $Y=0.1350 $X2=0.8370 $Y2=0.1350
r58 1 35 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8370 $Y=0.1350
+ $X2=0.8370 $Y2=0.1360
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.00420331f
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.00435743f
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%CLK VSS 10 3 8 5 1 6 7 4
c1 1 VSS 0.00255147f
c2 3 VSS 0.0597275f
c3 4 VSS 0.000976381f
c4 5 VSS 0.00409418f
c5 6 VSS 0.0040158f
c6 7 VSS 0.00226638f
c7 8 VSS 0.00210403f
r1 6 18 3.22357 $w=2.26279e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.2125 $X2=0.1080 $Y2=0.1820
r2 5 16 3.22357 $w=2.26279e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0575 $X2=0.1080 $Y2=0.0880
r3 17 18 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.1820 $X2=0.1080 $Y2=0.1820
r4 8 14 0.54189 $w=3.37e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1820 $X2=0.0810 $Y2=0.1630
r5 8 17 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1820 $X2=0.0945 $Y2=0.1820
r6 15 16 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.0880 $X2=0.1080 $Y2=0.0880
r7 7 15 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0880 $X2=0.0945 $Y2=0.0880
r8 13 14 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1530 $X2=0.0810 $Y2=0.1630
r9 12 13 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1530
r10 11 12 2.85657 $w=1.3e-08 $l=1.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1227 $X2=0.0810 $Y2=0.1350
r11 10 11 0.874462 $w=1.3e-08 $l=3.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1227
r12 10 4 1.57403 $w=1.3e-08 $l=6.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1122
r13 4 7 1.76614 $w=2.65738e-08 $l=2.42e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1122 $X2=0.0810 $Y2=0.0880
r14 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r15 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%PD2 VSS 7 12 4 1 5
c1 1 VSS 0.00724415f
c2 4 VSS 0.00187762f
c3 5 VSS 0.00234404f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4880 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r3 9 5 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.4605
+ $Y=0.2295 $X2=0.4860 $Y2=0.2295
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.4455
+ $Y=0.2295 $X2=0.4605 $Y2=0.2295
r5 1 8 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4320
+ $Y=0.2295 $X2=0.4455 $Y2=0.2295
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2295 $X2=0.4300 $Y2=0.2295
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2295 $X2=0.4175 $Y2=0.2295
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%MS VSS 10 41 44 49 51 13 17 18 14 3 15 12 1 4 11
+ 16
c1 1 VSS 0.0022044f
c2 3 VSS 0.00564576f
c3 4 VSS 0.00936411f
c4 10 VSS 0.0375471f
c5 11 VSS 0.00289897f
c6 12 VSS 0.00273297f
c7 13 VSS 0.00227538f
c8 14 VSS 0.00190588f
c9 15 VSS 0.00423695f
c10 16 VSS 0.00186513f
c11 17 VSS 0.00114364f
c12 18 VSS 0.000419751f
c13 19 VSS 0.00249555f
r1 51 50 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.2295 $X2=0.6625 $Y2=0.2295
r2 13 50 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6500 $Y=0.2295 $X2=0.6625 $Y2=0.2295
r3 12 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2295 $X2=0.5920 $Y2=0.2295
r4 49 12 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.2295 $X2=0.5795 $Y2=0.2295
r5 46 13 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6210 $Y=0.2295 $X2=0.6480 $Y2=0.2295
r6 4 46 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08 $X=0.5940
+ $Y=0.2295 $X2=0.6210 $Y2=0.2295
r7 4 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2295
+ $X2=0.5965 $Y2=0.2340
r8 15 19 4.48182 $w=1.47708e-08 $l=2.45051e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5965 $Y=0.2340 $X2=0.6210 $Y2=0.2335
r9 44 43 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.0405 $X2=0.6085 $Y2=0.0405
r10 42 43 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6040 $Y=0.0405 $X2=0.6085 $Y2=0.0405
r11 3 42 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5920 $Y=0.0405 $X2=0.6040 $Y2=0.0405
r12 11 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.0405 $X2=0.5920 $Y2=0.0405
r13 41 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0405 $X2=0.5795 $Y2=0.0405
r14 19 36 0.983973 $w=1.77222e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.2335 $X2=0.6210 $Y2=0.2245
r15 3 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0405
+ $X2=0.5940 $Y2=0.0540
r16 35 36 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.2135 $X2=0.6210 $Y2=0.2245
r17 34 35 6.64591 $w=1.3e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1850 $X2=0.6210 $Y2=0.2135
r18 33 34 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1660 $X2=0.6210 $Y2=0.1850
r19 32 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1525 $X2=0.6210 $Y2=0.1660
r20 31 32 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1310 $X2=0.6210 $Y2=0.1525
r21 30 31 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1115 $X2=0.6210 $Y2=0.1310
r22 17 28 1.15159 $w=1.75e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1000 $X2=0.6210 $Y2=0.0900
r23 17 30 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1000 $X2=0.6210 $Y2=0.1115
r24 16 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0540 $X2=0.5940 $Y2=0.0720
r25 27 28 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6075 $Y=0.0900 $X2=0.6210 $Y2=0.0900
r26 18 26 1.38478 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5940 $Y=0.0900 $X2=0.5830 $Y2=0.0900
r27 18 27 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5940 $Y=0.0900 $X2=0.6075 $Y2=0.0900
r28 18 29 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0900 $X2=0.5940 $Y2=0.0720
r29 25 26 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5515
+ $Y=0.0900 $X2=0.5830 $Y2=0.0900
r30 24 25 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0900 $X2=0.5515 $Y2=0.0900
r31 14 24 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5000
+ $Y=0.0900 $X2=0.5130 $Y2=0.0900
r32 1 21 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.5130
+ $Y=0.0900 $X2=0.5130 $Y2=0.0900
r33 1 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.0900
+ $X2=0.5130 $Y2=0.0900
r34 10 21 0.314665 $w=2.27e-07 $l=4.5e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5130 $Y2=0.0900
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%PD1 VSS 7 10 5 4 1
c1 1 VSS 0.0105868f
c2 4 VSS 0.00318439f
c3 5 VSS 0.00186088f
r1 10 9 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r2 8 9 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r3 5 8 0.123457 $w=8.1e-08 $l=1e-08 $layer=N_src_drn $thickness=1e-09 $X=0.3780
+ $Y=0.0675 $X2=0.3880 $Y2=0.0675
r4 4 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3220 $Y2=0.0675
r5 7 4 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r6 1 5 1e-05
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%MH VSS 9 50 54 60 64 10 18 14 12 3 4 15 16 19 17
+ 20 1
c1 1 VSS 0.000371526f
c2 3 VSS 0.00570406f
c3 4 VSS 0.00539951f
c4 9 VSS 0.0364537f
c5 10 VSS 0.00226024f
c6 11 VSS 8.96572e-20
c7 12 VSS 0.00279153f
c8 13 VSS 6.86277e-20
c9 14 VSS 0.00739289f
c10 15 VSS 0.00140629f
c11 16 VSS 0.000681003f
c12 17 VSS 0.000553846f
c13 18 VSS 0.00614736f
c14 19 VSS 2.3044e-20
c15 20 VSS 0.00289734f
r1 64 63 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r2 62 63 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r3 3 62 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3760 $Y=0.2295 $X2=0.3880 $Y2=0.2295
r4 13 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2295 $X2=0.3760 $Y2=0.2295
r5 58 59 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r6 60 58 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.1890 $X2=0.3635 $Y2=0.1890
r7 12 59 0.185185 $w=5.4e-08 $l=1e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r8 12 3 0.518519 $w=3.9e-08 $l=4.05494e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.1890 $X2=0.3760 $Y2=0.2295
r9 3 46 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2295
+ $X2=0.3780 $Y2=0.2340
r10 54 53 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r11 52 53 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4420 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r12 4 52 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4300 $Y=0.0405 $X2=0.4420 $Y2=0.0405
r13 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0405 $X2=0.4300 $Y2=0.0405
r14 10 4 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0810 $X2=0.4300 $Y2=0.0810
r15 50 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0810 $X2=0.4175 $Y2=0.0810
r16 46 47 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r17 44 47 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r18 43 44 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4160
+ $Y=0.2340 $X2=0.4050 $Y2=0.2340
r19 14 20 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4340
+ $Y=0.2340 $X2=0.4590 $Y2=0.2340
r20 14 43 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4340
+ $Y=0.2340 $X2=0.4160 $Y2=0.2340
r21 4 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0405
+ $X2=0.4320 $Y2=0.0360
r22 20 35 3.01468 $w=1.741e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4590 $Y2=0.2140
r23 37 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4455 $Y2=0.0360
r24 18 32 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4590 $Y2=0.0630
r25 18 38 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4455 $Y2=0.0360
r26 34 35 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1850 $X2=0.4590 $Y2=0.2140
r27 33 34 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1660 $X2=0.4590 $Y2=0.1850
r28 16 19 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1525 $X2=0.4590 $Y2=0.1310
r29 16 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1525 $X2=0.4590 $Y2=0.1660
r30 31 32 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0900 $X2=0.4590 $Y2=0.0630
r31 30 31 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1025 $X2=0.4590 $Y2=0.0900
r32 15 19 2.78392 $w=1.56471e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1140 $X2=0.4590 $Y2=0.1310
r33 15 30 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1140 $X2=0.4590 $Y2=0.1025
r34 19 28 4.18306 $w=1.49565e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1310 $X2=0.4820 $Y2=0.1310
r35 27 28 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5000
+ $Y=0.1310 $X2=0.4820 $Y2=0.1310
r36 26 27 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1310 $X2=0.5000 $Y2=0.1310
r37 17 25 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1310 $X2=0.5670 $Y2=0.1310
r38 17 26 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1310 $X2=0.5130 $Y2=0.1310
r39 1 22 2.36633 $w=2.3e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.5670
+ $Y=0.1305 $X2=0.5670 $Y2=0.1305
r40 1 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1305
+ $X2=0.5670 $Y2=0.1310
r41 9 22 0.314665 $w=2.27e-07 $l=4.5e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5670 $Y=0.1350 $X2=0.5670 $Y2=0.1305
r42 3 12 1e-05
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%CLKN VSS 13 14 15 77 79 8 22 26 7 17 1 16 19 20
+ 21 18 28 23 2 24 3
c1 1 VSS 0.00160348f
c2 2 VSS 6.0473e-20
c3 3 VSS 0.000170899f
c4 7 VSS 0.00756747f
c5 8 VSS 0.00787332f
c6 13 VSS 0.0597498f
c7 14 VSS 0.00440212f
c8 15 VSS 0.00458593f
c9 16 VSS 0.00585435f
c10 17 VSS 0.00577701f
c11 18 VSS 0.00522554f
c12 19 VSS 0.00342087f
c13 20 VSS 0.00448003f
c14 21 VSS 0.00455887f
c15 22 VSS 0.000598971f
c16 23 VSS 0.000578762f
c17 24 VSS 0.00143082f
c18 25 VSS 0.00351911f
c19 26 VSS 0.00152377f
c20 27 VSS 0.00374398f
c21 28 VSS 0.0230073f
r1 79 78 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r2 17 78 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r3 77 76 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r4 16 76 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r5 8 74 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0550 $Y2=0.2340
r6 7 71 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0550 $Y2=0.0360
r7 73 74 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.2340 $X2=0.0550 $Y2=0.2340
r8 21 73 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0460 $Y2=0.2340
r9 21 27 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0180 $Y2=0.2340
r10 70 71 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.0360 $X2=0.0550 $Y2=0.0360
r11 20 70 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0460 $Y2=0.0360
r12 20 25 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0180 $Y2=0.0360
r13 27 63 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.2340 $X2=0.0180 $Y2=0.2125
r14 25 61 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.0360 $X2=0.0180 $Y2=0.0575
r15 3 58 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6750 $Y=0.1350
+ $X2=0.6750 $Y2=0.1440
r16 15 3 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6750
+ $Y=0.1350 $X2=0.6750 $Y2=0.1350
r17 2 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
r18 14 2 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r19 62 63 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1820 $X2=0.0180 $Y2=0.2125
r20 19 26 0.998523 $w=1.74118e-08 $l=1.01119e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1630 $X2=0.0165 $Y2=0.1530
r21 19 62 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1630 $X2=0.0180 $Y2=0.1820
r22 60 61 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0880 $X2=0.0180 $Y2=0.0575
r23 18 26 5.19594 $w=1.44151e-08 $l=2.80401e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1250 $X2=0.0165 $Y2=0.1530
r24 18 60 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1250 $X2=0.0180 $Y2=0.0880
r25 24 58 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1135 $X2=0.6750 $Y2=0.1440
r26 23 56 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1530
r27 52 53 1.90199 $w=1.38333e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.0255 $Y=0.1530 $X2=0.0345 $Y2=0.1530
r28 26 52 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0165
+ $Y=0.1530 $X2=0.0255 $Y2=0.1530
r29 50 58 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.6750 $Y=0.1530
+ $X2=0.6750 $Y2=0.1440
r30 49 50 18.3054 $w=1.3e-08 $l=7.85e-08 $layer=M2 $thickness=3.6e-08 $X=0.5965
+ $Y=0.1530 $X2=0.6750 $Y2=0.1530
r31 48 49 29.3819 $w=1.3e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.4705
+ $Y=0.1530 $X2=0.5965 $Y2=0.1530
r32 47 48 15.2739 $w=1.3e-08 $l=6.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1530 $X2=0.4705 $Y2=0.1530
r33 47 56 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4050 $Y=0.1530
+ $X2=0.4050 $Y2=0.1530
r34 46 47 27.8662 $w=1.3e-08 $l=1.195e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.2855 $Y=0.1530 $X2=0.4050 $Y2=0.1530
r35 45 46 27.5164 $w=1.3e-08 $l=1.18e-07 $layer=M2 $thickness=3.6e-08 $X=0.1675
+ $Y=0.1530 $X2=0.2855 $Y2=0.1530
r36 44 45 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M2 $thickness=3.6e-08 $X=0.1510
+ $Y=0.1530 $X2=0.1675 $Y2=0.1530
r37 43 44 13.7582 $w=1.3e-08 $l=5.9e-08 $layer=M2 $thickness=3.6e-08 $X=0.0920
+ $Y=0.1530 $X2=0.1510 $Y2=0.1530
r38 42 43 13.7582 $w=1.3e-08 $l=5.9e-08 $layer=M2 $thickness=3.6e-08 $X=0.0330
+ $Y=0.1530 $X2=0.0920 $Y2=0.1530
r39 42 53 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.0330 $Y=0.1530
+ $X2=0.0345 $Y2=0.1530
r40 28 42 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.0215
+ $Y=0.1530 $X2=0.0330 $Y2=0.1530
r41 39 44 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1510 $Y=0.1440
+ $X2=0.1510 $Y2=0.1530
r42 22 39 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1510
+ $Y=0.1160 $X2=0.1510 $Y2=0.1440
r43 37 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1550 $Y=0.1350
+ $X2=0.1510 $Y2=0.1440
r44 36 37 4.43042 $w=1.53e-08 $l=7.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1475 $Y=0.1350 $X2=0.1550 $Y2=0.1350
r45 34 36 1.86855 $w=1.78125e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1435 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r46 1 34 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.1335
+ $Y=0.1350 $X2=0.1435 $Y2=0.1350
r47 13 1 2.53453 $w=1.32811e-07 $l=1.5e-09 $layer=LIG $thickness=5.23243e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1335 $Y2=0.1350
r48 13 36 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r49 8 17 1e-05
r50 7 16 1e-05
.ends

.subckt PM_DFFHQx4_ASAP7_75t_R%CLKB VSS 14 15 16 17 81 83 18 20 26 6 7 23 24 4
+ 25 22 19 1 21 2 8
c1 1 VSS 0.00174874f
c2 2 VSS 0.000781811f
c3 3 VSS 0.000732856f
c4 4 VSS 0.00115406f
c5 6 VSS 0.00861686f
c6 7 VSS 0.00863605f
c7 8 VSS 0.00501995f
c8 14 VSS 0.00601741f
c9 15 VSS 0.00582016f
c10 16 VSS 0.00507622f
c11 17 VSS 0.00591658f
c12 18 VSS 0.00542334f
c13 19 VSS 0.00542085f
c14 20 VSS 0.00399833f
c15 21 VSS 0.00331054f
c16 22 VSS 0.00278046f
c17 23 VSS 0.00745054f
c18 24 VSS 0.00560159f
c19 25 VSS 0.00125264f
c20 26 VSS 0.00546606f
r1 19 7 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1600 $Y2=0.2160
r2 83 19 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r3 18 6 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1600 $Y2=0.0540
r4 81 18 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r5 4 79 2.78395 $w=2.4e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08 $X=0.7290
+ $Y=0.1780 $X2=0.7250 $Y2=0.1780
r6 17 4 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.7290 $Y=0.1350 $X2=0.7290 $Y2=0.1780
r7 3 72 10.3807 $w=2.30357e-08 $l=0 $layer=LISD $thickness=3.675e-08 $X=0.6210
+ $Y=0.1780 $X2=0.6210 $Y2=0.1780
r8 16 3 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.6210 $Y=0.1350 $X2=0.6210 $Y2=0.1780
r9 2 65 2.78395 $w=2.4e-08 $l=5e-09 $layer=LIG $thickness=4.8e-08 $X=0.4590
+ $Y=0.1780 $X2=0.4640 $Y2=0.1780
r10 15 2 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4590 $Y2=0.1780
r11 7 57 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1655 $Y2=0.2340
r12 6 53 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1655 $Y2=0.0360
r13 78 79 4.8113 $w=2.22e-08 $l=1.5e-09 $layer=LISD $thickness=2.7e-08
+ $X=0.7235 $Y=0.1780 $X2=0.7250 $Y2=0.1780
r14 77 78 10.8887 $w=2.22e-08 $l=2.15e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7020 $Y=0.1780 $X2=0.7235 $Y2=0.1780
r15 76 77 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6885 $Y=0.1780 $X2=0.7020 $Y2=0.1780
r16 75 76 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6750 $Y=0.1780 $X2=0.6885 $Y2=0.1780
r17 74 75 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6615 $Y=0.1780 $X2=0.6750 $Y2=0.1780
r18 73 74 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6480 $Y=0.1780 $X2=0.6615 $Y2=0.1780
r19 72 73 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6210 $Y=0.1780 $X2=0.6480 $Y2=0.1780
r20 71 72 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5940 $Y=0.1780 $X2=0.6210 $Y2=0.1780
r21 70 71 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5805 $Y=0.1780 $X2=0.5940 $Y2=0.1780
r22 69 70 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5670 $Y=0.1780 $X2=0.5805 $Y2=0.1780
r23 68 69 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5535 $Y=0.1780 $X2=0.5670 $Y2=0.1780
r24 67 68 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5400 $Y=0.1780 $X2=0.5535 $Y2=0.1780
r25 66 67 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5265 $Y=0.1780 $X2=0.5400 $Y2=0.1780
r26 64 65 10.3823 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4775 $Y=0.1780 $X2=0.4640 $Y2=0.1780
r27 63 64 11.142 $w=2.22e-08 $l=2.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4995 $Y=0.1780 $X2=0.4775 $Y2=0.1780
r28 62 66 1.51936 $w=2.22e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.5235
+ $Y=0.1780 $X2=0.5265 $Y2=0.1780
r29 61 62 5.31775 $w=2.22e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5130 $Y=0.1780 $X2=0.5235 $Y2=0.1780
r30 8 61 5.31775 $w=2.22e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5025 $Y=0.1780 $X2=0.5130 $Y2=0.1780
r31 8 63 1.51936 $w=2.22e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.5025
+ $Y=0.1780 $X2=0.4995 $Y2=0.1780
r32 57 58 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1655
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r33 24 50 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2340 $X2=0.1890 $Y2=0.2125
r34 24 58 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2340 $X2=0.1755 $Y2=0.2340
r35 53 54 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1655
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r36 23 49 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1890 $Y2=0.0575
r37 23 54 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1755 $Y2=0.0360
r38 51 61 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5130 $Y=0.1845
+ $X2=0.5130 $Y2=0.1780
r39 22 51 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1680 $X2=0.5130 $Y2=0.1845
r40 48 49 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0880 $X2=0.1890 $Y2=0.0575
r41 47 48 11.3097 $w=1.3e-08 $l=4.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1365 $X2=0.1890 $Y2=0.0880
r42 46 50 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1990 $X2=0.1890 $Y2=0.2125
r43 45 46 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1890 $X2=0.1890 $Y2=0.1990
r44 20 45 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1735 $X2=0.1890 $Y2=0.1890
r45 20 47 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1735 $X2=0.1890 $Y2=0.1365
r46 43 51 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.5130 $Y=0.1890
+ $X2=0.5130 $Y2=0.1845
r47 42 43 22.0364 $w=1.3e-08 $l=9.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.4185
+ $Y=0.1890 $X2=0.5130 $Y2=0.1890
r48 41 42 22.0364 $w=1.3e-08 $l=9.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1890 $X2=0.4185 $Y2=0.1890
r49 40 41 15.7403 $w=1.3e-08 $l=6.75e-08 $layer=M2 $thickness=3.6e-08 $X=0.2565
+ $Y=0.1890 $X2=0.3240 $Y2=0.1890
r50 39 40 15.7403 $w=1.3e-08 $l=6.75e-08 $layer=M2 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1890 $X2=0.2565 $Y2=0.1890
r51 39 45 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1890 $Y=0.1890
+ $X2=0.1890 $Y2=0.1890
r52 26 39 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.1775
+ $Y=0.1890 $X2=0.1890 $Y2=0.1890
r53 37 41 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.3240 $Y=0.1890
+ $X2=0.3240 $Y2=0.1890
r54 36 37 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1735 $X2=0.3240 $Y2=0.1890
r55 21 34 3.60008 $w=1.51951e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3240 $Y=0.1555 $X2=0.3240 $Y2=0.1350
r56 21 36 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1555 $X2=0.3240 $Y2=0.1735
r57 25 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r58 25 34 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3375 $Y=0.1350 $X2=0.3240 $Y2=0.1350
r59 14 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r60 1 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
.ends


*
.SUBCKT DFFHQx4_ASAP7_75t_R VSS VDD CLK D Q
*
* VSS VSS
* VDD VDD
* CLK CLK
* D D
* Q Q
*
*

MM20 N_MM20_d N_MM20_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM23 N_MM23_d N_MM22_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM10_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM6 N_MM6_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM12 N_MM12_d N_MM12_g N_MM12_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM17 N_MM17_d N_MM13_g N_MM17_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM16 N_MM16_d N_MM19_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM14 N_MM14_d N_MM14_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM24 N_MM24_d N_MM24_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@2 N_MM24@2_d N_MM24@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM38 N_MM38_d N_MM38_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM38@4 N_MM38@4_d N_MM38@4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM38@3 N_MM38@3_d N_MM38@3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM38@2 N_MM38@2_d N_MM38@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM21 N_MM21_d N_MM20_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM22 N_MM22_d N_MM22_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM13 N_MM13_d N_MM13_g N_MM13_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM18 N_MM18_d N_MM18_g N_MM18_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM19 N_MM19_d N_MM19_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM15 N_MM15_d N_MM14_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM25 N_MM25_d N_MM24_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@2 N_MM25@2_d N_MM24@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM37 N_MM37_d N_MM38_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM37@4 N_MM37@4_d N_MM38@4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM37@3 N_MM37@3_d N_MM38@3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM37@2 N_MM37@2_d N_MM38@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "DFFHQx4_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "DFFHQx4_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_DFFHQx4_ASAP7_75t_R%noxref_29 VSS N_noxref_29_1
+ PM_DFFHQx4_ASAP7_75t_R%noxref_29
cc_1 N_noxref_29_1 N_MM38@2_g 0.00146974f
cc_2 N_noxref_29_1 N_Q_14 0.000820897f
x_PM_DFFHQx4_ASAP7_75t_R%noxref_30 VSS N_noxref_30_1
+ PM_DFFHQx4_ASAP7_75t_R%noxref_30
cc_3 N_noxref_30_1 N_MM38@2_g 0.00147125f
cc_4 N_noxref_30_1 N_Q_16 0.000827693f
cc_5 N_noxref_30_1 N_noxref_29_1 0.00176533f
x_PM_DFFHQx4_ASAP7_75t_R%Q VSS Q N_MM38_d N_MM38@4_d N_MM38@3_d N_MM38@2_d
+ N_MM37@3_d N_MM37@2_d N_MM37_d N_MM37@4_d N_Q_14 N_Q_18 N_Q_16 N_Q_15 N_Q_13
+ N_Q_21 N_Q_20 N_Q_2 N_Q_3 N_Q_4 N_Q_1 PM_DFFHQx4_ASAP7_75t_R%Q
cc_6 N_Q_14 N_NET049_1 0.000617828f
cc_7 N_Q_18 N_MM38@3_g 0.000637856f
cc_8 N_Q_16 N_MM38@3_g 0.0305284f
cc_9 N_Q_15 N_MM38_g 0.0306721f
cc_10 N_Q_13 N_MM38_g 0.0672423f
cc_11 N_Q_21 N_NET049_22 0.00105729f
cc_12 N_Q_20 N_NET049_20 0.00107366f
cc_13 N_Q_2 N_NET049_19 0.0016909f
cc_14 N_Q_3 N_MM38@3_g 0.00183993f
cc_15 N_Q_4 N_MM38@3_g 0.0019328f
cc_16 N_Q_1 N_MM38_g 0.00222651f
cc_17 N_Q_2 N_MM38_g 0.00231374f
cc_18 N_Q_21 N_NET049_18 0.00247279f
cc_19 N_Q_20 N_NET049_17 0.00258362f
cc_20 N_Q_16 N_NET049_1 0.00958051f
cc_21 N_Q_14 N_MM38@2_g 0.0367693f
cc_22 N_Q_13 N_MM38@4_g 0.0367935f
cc_23 N_Q_14 N_MM38@3_g 0.0700176f
x_PM_DFFHQx4_ASAP7_75t_R%PD3 VSS N_MM9_s N_MM8_d N_PD3_1
+ PM_DFFHQx4_ASAP7_75t_R%PD3
cc_24 N_PD3_1 N_MM9_g 0.00776936f
cc_25 N_PD3_1 N_MM11_g 0.00769417f
x_PM_DFFHQx4_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_DFFHQx4_ASAP7_75t_R%noxref_23
cc_26 N_noxref_23_1 N_MM3_g 0.00183986f
cc_27 N_noxref_23_1 N_CLKB_6 0.000100385f
cc_28 N_noxref_23_1 N_CLKB_18 0.000557096f
cc_29 N_noxref_23_1 N_noxref_21_1 0.0076962f
cc_30 N_noxref_23_1 N_noxref_22_1 0.000463105f
x_PM_DFFHQx4_ASAP7_75t_R%PD4 VSS N_MM18_s N_MM19_d N_PD4_1
+ PM_DFFHQx4_ASAP7_75t_R%PD4
cc_31 N_PD4_1 N_MM18_g 0.00777916f
cc_32 N_PD4_1 N_MM19_g 0.00770946f
x_PM_DFFHQx4_ASAP7_75t_R%PU1 VSS N_MM3_d N_MM1_s N_PU1_1
+ PM_DFFHQx4_ASAP7_75t_R%PU1
cc_33 N_PU1_1 N_MM3_g 0.0172559f
cc_34 N_PU1_1 N_MM1_g 0.0169761f
x_PM_DFFHQx4_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_DFFHQx4_ASAP7_75t_R%noxref_24
cc_35 N_noxref_24_1 N_MM3_g 0.00185815f
cc_36 N_noxref_24_1 N_CLKB_7 0.000106992f
cc_37 N_noxref_24_1 N_CLKB_19 0.000554117f
cc_38 N_noxref_24_1 N_noxref_21_1 0.000462747f
cc_39 N_noxref_24_1 N_noxref_22_1 0.00769003f
cc_40 N_noxref_24_1 N_noxref_23_1 0.00121513f
x_PM_DFFHQx4_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_DFFHQx4_ASAP7_75t_R%noxref_21
cc_41 N_noxref_21_1 N_CLKN_1 0.000375521f
cc_42 N_noxref_21_1 N_MM22_g 0.00344449f
cc_43 N_noxref_21_1 N_CLKB_6 0.000343025f
cc_44 N_noxref_21_1 N_CLKB_18 0.0270493f
x_PM_DFFHQx4_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_DFFHQx4_ASAP7_75t_R%noxref_22
cc_45 N_noxref_22_1 N_CLKN_1 0.000376956f
cc_46 N_noxref_22_1 N_MM22_g 0.00344531f
cc_47 N_noxref_22_1 N_CLKB_7 0.000338042f
cc_48 N_noxref_22_1 N_CLKB_19 0.0270518f
cc_49 N_noxref_22_1 N_noxref_21_1 0.00143019f
x_PM_DFFHQx4_ASAP7_75t_R%D VSS D N_MM3_g N_D_5 N_D_6 N_D_7 N_D_9 N_D_1 N_D_4
+ N_D_8 PM_DFFHQx4_ASAP7_75t_R%D
cc_50 N_D_5 N_MM10_g 6.17104e-20
cc_51 N_D_5 N_CLKN_22 0.0001457f
cc_52 N_D_5 N_CLKN_23 7.16963e-20
cc_53 N_D_5 N_CLKN_1 0.000113233f
cc_54 N_D_6 N_CLKN_28 0.000662514f
cc_55 N_D_5 N_CLKN_28 0.00319312f
x_PM_DFFHQx4_ASAP7_75t_R%noxref_26 VSS N_noxref_26_1
+ PM_DFFHQx4_ASAP7_75t_R%noxref_26
cc_56 N_noxref_26_1 N_SS_11 0.0169261f
cc_57 N_noxref_26_1 N_SH_1 0.000201572f
cc_58 N_noxref_26_1 N_MM14_g 0.00603272f
cc_59 N_noxref_26_1 N_noxref_25_1 0.00154151f
x_PM_DFFHQx4_ASAP7_75t_R%noxref_28 VSS N_noxref_28_1
+ PM_DFFHQx4_ASAP7_75t_R%noxref_28
cc_60 N_noxref_28_1 N_SS_11 0.000654239f
cc_61 N_noxref_28_1 N_MM24_g 0.00171599f
cc_62 N_noxref_28_1 N_noxref_25_1 0.00047705f
cc_63 N_noxref_28_1 N_noxref_26_1 0.00776988f
cc_64 N_noxref_28_1 N_noxref_27_1 0.00123538f
x_PM_DFFHQx4_ASAP7_75t_R%noxref_27 VSS N_noxref_27_1
+ PM_DFFHQx4_ASAP7_75t_R%noxref_27
cc_65 N_noxref_27_1 N_SS_10 0.000649634f
cc_66 N_noxref_27_1 N_MM24_g 0.00170937f
cc_67 N_noxref_27_1 N_noxref_25_1 0.00777796f
cc_68 N_noxref_27_1 N_noxref_26_1 0.000481328f
x_PM_DFFHQx4_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_DFFHQx4_ASAP7_75t_R%noxref_25
cc_69 N_noxref_25_1 N_SS_10 0.0170399f
cc_70 N_noxref_25_1 N_MM14_g 0.00613146f
x_PM_DFFHQx4_ASAP7_75t_R%SS VSS N_MM19_g N_MM14_d N_MM15_d N_SS_10 N_SS_11
+ N_SS_4 N_SS_15 N_SS_3 N_SS_14 N_SS_1 N_SS_16 N_SS_12 N_SS_13
+ PM_DFFHQx4_ASAP7_75t_R%SS
cc_71 N_MM19_g N_CLKB_8 0.000226513f
cc_72 N_MM19_g N_CLKB_4 0.000532742f
cc_73 N_MM19_g N_MM18_g 0.0135372f
x_PM_DFFHQx4_ASAP7_75t_R%PD5 VSS N_MM17_s N_MM16_d N_PD5_4 N_PD5_1 N_PD5_5
+ PM_DFFHQx4_ASAP7_75t_R%PD5
cc_74 N_PD5_4 N_MM13_g 0.0152265f
cc_75 N_PD5_1 N_MM18_g 0.0006494f
cc_76 N_PD5_5 N_MM18_g 0.00692166f
cc_77 N_PD5_4 N_MM18_g 0.0239536f
cc_78 N_PD5_1 N_MM19_g 0.000890818f
cc_79 N_PD5_5 N_MM19_g 0.0156069f
cc_80 N_PD5_1 N_SH_14 0.000316294f
cc_81 N_PD5_1 N_SH_16 0.000448266f
cc_82 N_PD5_1 N_SH_17 0.000570122f
cc_83 N_PD5_4 N_SH_5 0.000659814f
cc_84 N_PD5_1 N_SH_25 0.00255748f
x_PM_DFFHQx4_ASAP7_75t_R%NET049 VSS N_MM38_g N_MM38@4_g N_MM38@3_g N_MM38@2_g
+ N_MM24_d N_MM24@2_d N_MM25_d N_MM25@2_d N_NET049_13 N_NET049_16 N_NET049_4
+ N_NET049_17 N_NET049_18 N_NET049_14 N_NET049_3 N_NET049_1 N_NET049_22
+ N_NET049_20 N_NET049_19 PM_DFFHQx4_ASAP7_75t_R%NET049
cc_85 N_NET049_13 N_SH_2 0.000390645f
cc_86 N_NET049_13 N_SH_23 0.000639185f
cc_87 N_NET049_13 N_MM24@2_g 0.0400009f
cc_88 N_NET049_16 N_SH_23 0.000498905f
cc_89 N_NET049_4 N_SH_2 0.000525096f
cc_90 N_NET049_17 N_SH_2 0.00054745f
cc_91 N_NET049_18 N_SH_2 0.000605994f
cc_92 N_NET049_16 N_SH_29 0.000746966f
cc_93 N_NET049_14 N_MM24_g 0.031445f
cc_94 N_NET049_4 N_SH_23 0.00112025f
cc_95 N_MM38_g N_MM24@2_g 0.0016573f
cc_96 N_NET049_3 N_MM24_g 0.0019584f
cc_97 N_NET049_4 N_MM24_g 0.00211694f
cc_98 N_NET049_14 N_SH_2 0.00514814f
cc_99 N_NET049_13 N_MM24_g 0.0697409f
x_PM_DFFHQx4_ASAP7_75t_R%SH VSS N_MM14_g N_MM24_g N_MM24@2_g N_MM13_s N_MM18_d
+ N_MM12_s N_MM17_d N_SH_5 N_SH_6 N_SH_19 N_SH_14 N_SH_15 N_SH_24 N_SH_26
+ N_SH_17 N_SH_18 N_SH_16 N_SH_22 N_SH_2 N_SH_28 N_SH_27 N_SH_21 N_SH_23 N_SH_1
+ N_SH_25 N_SH_20 N_SH_29 PM_DFFHQx4_ASAP7_75t_R%SH
cc_100 N_SH_5 N_CLKN_28 0.000133654f
cc_101 N_SH_6 N_MM13_g 0.000162566f
cc_102 N_SH_19 N_CLKN_24 0.00021084f
cc_103 N_SH_14 N_MM13_g 0.00676501f
cc_104 N_SH_15 N_MM13_g 0.00683707f
cc_105 N_SH_24 N_CLKN_24 0.000368027f
cc_106 N_SH_26 N_CLKN_24 0.000943177f
cc_107 N_SH_17 N_CLKN_3 0.000462074f
cc_108 N_SH_5 N_CLKN_3 0.000507775f
cc_109 N_SH_18 N_CLKN_24 0.000526869f
cc_110 N_SH_16 N_CLKN_24 0.000536657f
cc_111 N_SH_16 N_CLKN_28 0.00107497f
cc_112 N_SH_17 N_CLKN_24 0.00385053f
cc_113 N_SH_5 N_MM13_g 0.0184214f
cc_114 N_SH_15 N_CLKB_26 8.05469e-20
cc_115 N_SH_24 N_CLKB_8 0.000189181f
cc_116 N_SH_26 N_CLKB_8 0.000202748f
cc_117 N_SH_14 N_MM12_g 0.00679975f
cc_118 N_SH_6 N_CLKB_8 0.00030691f
cc_119 N_SH_19 N_CLKB_4 0.000412756f
cc_120 N_SH_17 N_CLKB_8 0.000427812f
cc_121 N_SH_18 N_CLKB_8 0.000603914f
cc_122 N_SH_15 N_CLKB_4 0.000926173f
cc_123 N_SH_6 N_MM18_g 0.000993639f
cc_124 N_SH_15 N_CLKB_8 0.00227596f
cc_125 N_SH_5 N_MM12_g 0.00950991f
cc_126 N_SH_15 N_MM18_g 0.0161925f
cc_127 N_SH_17 N_MS_3 0.000115732f
cc_128 N_SH_24 N_MS_3 0.000121935f
cc_129 N_SH_15 N_MS_3 0.000436461f
cc_130 N_SH_6 N_MS_3 0.000223628f
cc_131 N_SH_14 N_MS_3 0.000463628f
cc_132 N_SH_24 N_MS_4 0.000306661f
cc_133 N_SH_6 N_MS_4 0.000415496f
cc_134 N_SH_16 N_MS_16 0.000475592f
cc_135 N_SH_15 N_MS_4 0.000586807f
cc_136 N_SH_24 N_MS_17 0.000636321f
cc_137 N_SH_16 N_MS_18 0.00157051f
cc_138 N_SH_5 N_MS_3 0.00367882f
cc_139 N_SH_18 N_MM19_g 0.00013191f
cc_140 N_SH_22 N_MM19_g 0.000149903f
cc_141 N_SH_2 N_MM19_g 0.000157237f
cc_142 N_SH_28 N_MM19_g 0.000158626f
cc_143 N_SH_27 N_MM19_g 0.000209489f
cc_144 N_MM14_g N_SS_10 0.00676633f
cc_145 N_MM14_g N_SS_11 0.00687495f
cc_146 N_SH_21 N_SS_4 0.000263418f
cc_147 N_SH_2 N_SS_15 0.000282312f
cc_148 N_SH_23 N_SS_15 0.00154407f
cc_149 N_SH_22 N_SS_15 0.00675605f
cc_150 N_MM14_g N_SS_3 0.000398578f
cc_151 N_MM14_g N_SS_4 0.000500791f
cc_152 N_SH_21 N_SS_14 0.000659405f
cc_153 N_SH_1 N_SS_1 0.000680601f
cc_154 N_SH_25 N_SS_16 0.000802451f
cc_155 N_SH_17 N_SS_1 0.000843506f
cc_156 N_SH_28 N_SS_15 0.000908679f
cc_157 N_SH_20 N_SS_12 0.000963811f
cc_158 N_SH_20 N_SS_13 0.00099593f
cc_159 N_MM14_g N_SS_1 0.00117266f
cc_160 N_SH_1 N_MM19_g 0.00129033f
cc_161 N_SH_28 N_SS_14 0.00133106f
cc_162 N_SH_19 N_SS_12 0.00154575f
cc_163 N_SH_29 N_SS_15 0.001873f
cc_164 N_SH_17 N_SS_12 0.00488306f
cc_165 N_MM14_g N_MM19_g 0.0294575f
x_PM_DFFHQx4_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_DFFHQx4_ASAP7_75t_R%noxref_19
cc_166 N_noxref_19_1 N_MM20_g 0.00369121f
cc_167 N_noxref_19_1 N_CLKN_19 6.23838e-20
cc_168 N_noxref_19_1 N_CLKN_18 0.000314677f
cc_169 N_noxref_19_1 N_CLKN_7 0.000504056f
cc_170 N_noxref_19_1 N_CLKN_16 0.0277516f
x_PM_DFFHQx4_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_DFFHQx4_ASAP7_75t_R%noxref_20
cc_171 N_noxref_20_1 N_MM20_g 0.0036696f
cc_172 N_noxref_20_1 N_CLKN_26 8.90152e-20
cc_173 N_noxref_20_1 N_CLKN_18 0.000152903f
cc_174 N_noxref_20_1 N_CLKN_19 0.000197677f
cc_175 N_noxref_20_1 N_CLKN_8 0.000426905f
cc_176 N_noxref_20_1 N_CLKN_17 0.0276789f
cc_177 N_noxref_20_1 N_noxref_19_1 0.0020412f
x_PM_DFFHQx4_ASAP7_75t_R%CLK VSS CLK N_MM20_g N_CLK_8 N_CLK_5 N_CLK_1 N_CLK_6
+ N_CLK_7 N_CLK_4 PM_DFFHQx4_ASAP7_75t_R%CLK
x_PM_DFFHQx4_ASAP7_75t_R%PD2 VSS N_MM10_s N_MM11_d N_PD2_4 N_PD2_1 N_PD2_5
+ PM_DFFHQx4_ASAP7_75t_R%PD2
cc_178 N_PD2_4 N_MM10_g 0.0149608f
cc_179 N_PD2_4 N_CLKB_8 0.000148366f
cc_180 N_PD2_1 N_CLKB_2 0.00053908f
cc_181 N_PD2_5 N_CLKB_8 0.00129266f
cc_182 N_PD2_1 N_MM9_g 0.0020703f
cc_183 N_PD2_5 N_MM9_g 0.00736383f
cc_184 N_PD2_4 N_MM9_g 0.0238877f
cc_185 N_PD2_5 N_MM11_g 0.0147541f
cc_186 N_PD2_1 N_MH_14 0.000447355f
cc_187 N_PD2_4 N_MH_3 0.000608221f
cc_188 N_PD2_1 N_MH_20 0.00321259f
x_PM_DFFHQx4_ASAP7_75t_R%MS VSS N_MM11_g N_MM6_d N_MM12_d N_MM7_d N_MM13_d
+ N_MS_13 N_MS_17 N_MS_18 N_MS_14 N_MS_3 N_MS_15 N_MS_12 N_MS_1 N_MS_4 N_MS_11
+ N_MS_16 PM_DFFHQx4_ASAP7_75t_R%MS
cc_189 N_MS_13 N_CLKN_24 0.000300156f
cc_190 N_MS_13 N_MM10_g 0.000129709f
cc_191 N_MS_13 N_CLKN_3 0.000187441f
cc_192 N_MS_13 N_CLKN_28 0.000242052f
cc_193 N_MS_17 N_CLKN_3 0.000264376f
cc_194 N_MS_17 N_CLKN_24 0.00466327f
cc_195 N_MS_18 N_CLKN_24 0.000633343f
cc_196 N_MS_14 N_CLKN_28 0.0025845f
cc_197 N_MS_13 N_MM13_g 0.0155539f
cc_198 N_MS_3 N_CLKB_22 0.000224759f
cc_199 N_MS_3 N_CLKB_8 0.000486976f
cc_200 N_MS_3 N_CLKB_2 0.000122475f
cc_201 N_MS_3 N_MM9_g 0.000156839f
cc_202 N_MS_3 N_CLKB_26 0.000176268f
cc_203 N_MS_15 N_CLKB_22 0.000275574f
cc_204 N_MS_13 N_MM12_g 0.00788347f
cc_205 N_MS_12 N_MM12_g 0.00779128f
cc_206 N_MS_15 N_CLKB_8 0.000390917f
cc_207 N_MS_1 N_MM9_g 0.000565744f
cc_208 N_MS_17 N_CLKB_8 0.00156161f
cc_209 N_MS_4 N_MM12_g 0.00248674f
cc_210 N_MS_11 N_MM12_g 0.00651039f
cc_211 N_MS_4 N_CLKB_8 0.00634067f
cc_212 N_MM11_g N_MM9_g 0.0142124f
cc_213 N_MS_3 N_MM12_g 0.0259694f
x_PM_DFFHQx4_ASAP7_75t_R%PD1 VSS N_MM5_d N_MM4_s N_PD1_5 N_PD1_4 N_PD1_1
+ PM_DFFHQx4_ASAP7_75t_R%PD1
cc_214 N_PD1_5 N_CLKN_2 0.000865609f
cc_215 N_PD1_5 N_CLKN_23 0.000308608f
cc_216 N_PD1_5 N_MM10_g 0.0343911f
cc_217 N_PD1_4 N_D_1 0.00079009f
cc_218 N_PD1_4 N_MM3_g 0.0350575f
cc_219 N_PD1_4 N_CLKB_25 0.000422018f
cc_220 N_PD1_4 N_CLKB_1 0.002016f
cc_221 N_PD1_4 N_MM1_g 0.0737201f
cc_222 N_PD1_1 N_MH_4 0.00122819f
cc_223 N_PD1_1 N_MH_10 0.00350642f
x_PM_DFFHQx4_ASAP7_75t_R%MH VSS N_MM7_g N_MM4_d N_MM9_d N_MM1_d N_MM10_d
+ N_MH_10 N_MH_18 N_MH_14 N_MH_12 N_MH_3 N_MH_4 N_MH_15 N_MH_16 N_MH_19 N_MH_17
+ N_MH_20 N_MH_1 PM_DFFHQx4_ASAP7_75t_R%MH
cc_224 N_MH_10 N_CLKN_3 9.78342e-20
cc_225 N_MH_10 N_CLKN_28 0.000116793f
cc_226 N_MH_10 N_MM13_g 0.000161351f
cc_227 N_MH_10 N_CLKN_23 0.000329309f
cc_228 N_MH_18 N_CLKN_23 0.00034899f
cc_229 N_MH_14 N_CLKN_23 0.000411476f
cc_230 N_MH_12 N_MM10_g 0.0164399f
cc_231 N_MH_3 N_CLKN_2 0.000843464f
cc_232 N_MH_4 N_MM10_g 0.00108194f
cc_233 N_MH_15 N_CLKN_23 0.00117172f
cc_234 N_MH_3 N_MM10_g 0.00123791f
cc_235 N_MH_16 N_CLKN_23 0.00127743f
cc_236 N_MH_10 N_CLKN_2 0.00161224f
cc_237 N_MH_19 N_CLKN_23 0.0029272f
cc_238 N_MH_17 N_CLKN_28 0.00353864f
cc_239 N_MH_10 N_MM10_g 0.0529361f
cc_240 N_MH_10 N_CLKB_22 0.000382658f
cc_241 N_MH_10 N_CLKB_21 0.000148803f
cc_242 N_MH_10 N_MM1_g 0.000431753f
cc_243 N_MH_10 N_CLKB_25 0.000288941f
cc_244 N_MH_16 N_CLKB_22 0.0026235f
cc_245 N_MH_3 N_CLKB_1 0.000337537f
cc_246 N_MH_20 N_CLKB_22 0.000355692f
cc_247 N_MH_17 N_CLKB_8 0.000623313f
cc_248 N_MH_1 N_CLKB_8 0.00222084f
cc_249 N_MH_4 N_MM9_g 0.000631901f
cc_250 N_MH_3 N_CLKB_21 0.000654326f
cc_251 N_MH_12 N_CLKB_1 0.000792606f
cc_252 N_MH_16 N_CLKB_2 0.00079907f
cc_253 N_MH_3 N_MM1_g 0.00173126f
cc_254 N_MH_14 N_CLKB_26 0.00280554f
cc_255 N_MH_17 N_CLKB_22 0.00362113f
cc_256 N_MM7_g N_CLKB_8 0.00464795f
cc_257 N_MH_12 N_MM1_g 0.0337437f
cc_258 N_MM7_g N_MM12_g 0.0127649f
cc_259 N_MH_10 N_MM9_g 0.0364406f
cc_260 N_MH_4 N_MS_1 0.000395735f
cc_261 N_MH_17 N_MS_18 0.000495525f
cc_262 N_MH_17 N_MS_1 0.000817008f
cc_263 N_MM7_g N_MS_3 0.000858853f
cc_264 N_MH_1 N_MS_14 0.00102972f
cc_265 N_MH_17 N_MS_17 0.00103636f
cc_266 N_MH_1 N_MM11_g 0.00115617f
cc_267 N_MM7_g N_MS_1 0.00117893f
cc_268 N_MH_15 N_MS_14 0.00123415f
cc_269 N_MM7_g N_MS_12 0.00633402f
cc_270 N_MM7_g N_MS_11 0.00642325f
cc_271 N_MH_17 N_MS_14 0.00719832f
cc_272 N_MM7_g N_MM11_g 0.0294283f
x_PM_DFFHQx4_ASAP7_75t_R%CLKN VSS N_MM22_g N_MM10_g N_MM13_g N_MM20_d N_MM21_d
+ N_CLKN_8 N_CLKN_22 N_CLKN_26 N_CLKN_7 N_CLKN_17 N_CLKN_1 N_CLKN_16 N_CLKN_19
+ N_CLKN_20 N_CLKN_21 N_CLKN_18 N_CLKN_28 N_CLKN_23 N_CLKN_2 N_CLKN_24 N_CLKN_3
+ PM_DFFHQx4_ASAP7_75t_R%CLKN
cc_273 N_CLKN_8 N_MM20_g 0.00110864f
cc_274 N_CLKN_22 N_MM20_g 0.000245351f
cc_275 N_CLKN_26 N_MM20_g 0.000250533f
cc_276 N_CLKN_7 N_MM20_g 0.00112439f
cc_277 N_CLKN_17 N_MM20_g 0.0112181f
cc_278 N_CLKN_1 N_MM20_g 0.000334106f
cc_279 N_CLKN_16 N_MM20_g 0.011223f
cc_280 N_CLKN_19 N_CLK_8 0.000503194f
cc_281 N_CLKN_20 N_CLK_5 0.000802024f
cc_282 N_CLKN_26 N_CLK_1 0.000820681f
cc_283 N_CLKN_21 N_CLK_6 0.000823953f
cc_284 N_CLKN_21 N_CLK_8 0.000841621f
cc_285 N_CLKN_22 N_CLK_7 0.00105095f
cc_286 N_CLKN_18 N_CLK_7 0.00115986f
cc_287 N_CLKN_26 N_CLK_8 0.00159419f
cc_288 N_CLKN_28 N_CLK_8 0.00182173f
cc_289 N_CLKN_1 N_CLK_1 0.00252778f
cc_290 N_CLKN_20 N_CLK_7 0.00268911f
cc_291 N_CLKN_22 N_CLK_8 0.00310543f
cc_292 N_CLKN_26 N_CLK_4 0.00358108f
cc_293 N_MM22_g N_MM20_g 0.0350376f
x_PM_DFFHQx4_ASAP7_75t_R%CLKB VSS N_MM1_g N_MM9_g N_MM12_g N_MM18_g N_MM23_d
+ N_MM22_d N_CLKB_18 N_CLKB_20 N_CLKB_26 N_CLKB_6 N_CLKB_7 N_CLKB_23 N_CLKB_24
+ N_CLKB_4 N_CLKB_25 N_CLKB_22 N_CLKB_19 N_CLKB_1 N_CLKB_21 N_CLKB_2 N_CLKB_8
+ PM_DFFHQx4_ASAP7_75t_R%CLKB
cc_294 N_CLKB_18 N_CLK_6 8.57401e-20
cc_295 N_CLKB_20 N_CLK_6 8.70575e-20
cc_296 N_CLKB_26 N_CLK_6 0.000118898f
cc_297 N_CLKB_6 N_CLK_6 0.000381852f
cc_298 N_CLKB_7 N_CLK_6 0.000381549f
cc_299 N_CLKB_23 N_CLK_7 0.000503611f
cc_300 N_CLKB_20 N_CLK_8 0.000505036f
cc_301 N_CLKB_23 N_CLK_5 0.00118598f
cc_302 N_CLKB_24 N_CLK_6 0.00193195f
cc_303 N_CLKB_24 N_MM22_g 4.19348e-20
cc_304 N_CLKB_6 N_MM22_g 0.000752161f
cc_305 N_CLKB_7 N_MM22_g 0.000767599f
cc_306 N_CLKB_4 N_MM13_g 0.000219293f
cc_307 N_CLKB_25 N_CLKN_28 0.000266311f
cc_308 N_CLKB_22 N_CLKN_28 0.000670286f
cc_309 N_CLKB_24 N_CLKN_22 0.000319149f
cc_310 N_CLKB_23 N_CLKN_22 0.000357074f
cc_311 N_CLKB_19 N_MM22_g 0.0112354f
cc_312 N_CLKB_1 N_CLKN_2 0.00165233f
cc_313 N_CLKB_21 N_CLKN_28 0.0010429f
cc_314 N_CLKB_20 N_CLKN_22 0.00771889f
cc_315 N_CLKB_25 N_CLKN_2 0.000497806f
cc_316 N_CLKB_20 N_CLKN_28 0.000511038f
cc_317 N_CLKB_2 N_MM10_g 0.000569193f
cc_318 N_CLKB_8 N_CLKN_24 0.00057155f
cc_319 N_CLKB_8 N_CLKN_3 0.00269812f
cc_320 N_CLKB_26 N_CLKN_23 0.000627932f
cc_321 N_CLKB_20 N_CLKN_1 0.00087742f
cc_322 N_CLKB_19 N_CLKN_1 0.00109806f
cc_323 N_CLKB_25 N_CLKN_23 0.00264648f
cc_324 N_MM9_g N_MM10_g 0.00369689f
cc_325 N_CLKB_8 N_MM13_g 0.00422515f
cc_326 N_MM18_g N_MM13_g 0.00583568f
cc_327 N_MM1_g N_MM10_g 0.00703134f
cc_328 N_MM12_g N_MM13_g 0.0183392f
cc_329 N_CLKB_26 N_CLKN_28 0.0308884f
cc_330 N_CLKB_18 N_MM22_g 0.0389352f
cc_331 N_CLKB_21 N_MM3_g 0.000133069f
cc_332 N_CLKB_7 N_MM3_g 0.000140716f
cc_333 N_CLKB_20 N_MM3_g 0.000201121f
cc_334 N_CLKB_1 N_MM3_g 0.000269558f
cc_335 N_CLKB_25 N_MM3_g 0.000620612f
cc_336 N_CLKB_23 N_D_7 0.000918792f
cc_337 N_CLKB_26 N_D_6 0.00107356f
cc_338 N_CLKB_21 N_D_6 0.00114524f
cc_339 N_CLKB_24 N_D_9 0.00121775f
cc_340 N_CLKB_1 N_D_1 0.00161522f
cc_341 N_CLKB_20 N_D_4 0.00183283f
cc_342 N_CLKB_25 N_D_6 0.00202843f
cc_343 N_CLKB_20 N_D_5 0.00243182f
cc_344 N_CLKB_20 N_D_8 0.00403363f
cc_345 N_MM1_g N_MM3_g 0.00526968f
*END of DFFHQx4_ASAP7_75t_R.pxi
.ENDS
** Design:	DFFLQNx1_ASAP7_75t_R
* Created:	"Fri Aug 17 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "DFFLQNx1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "DFFLQNx1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_DFFLQNx1_ASAP7_75t_R%noxref_29 VSS 1
c1 1 VSS 0.00452565f
.ends

.subckt PM_DFFLQNx1_ASAP7_75t_R%noxref_28 VSS 1
c1 1 VSS 0.00477285f
.ends

.subckt PM_DFFLQNx1_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.041809f
.ends

.subckt PM_DFFLQNx1_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.041851f
.ends

.subckt PM_DFFLQNx1_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.00423879f
.ends

.subckt PM_DFFLQNx1_ASAP7_75t_R%noxref_26 VSS 1
c1 1 VSS 0.0415041f
.ends

.subckt PM_DFFLQNx1_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.00434691f
.ends

.subckt PM_DFFLQNx1_ASAP7_75t_R%noxref_27 VSS 1
c1 1 VSS 0.0415016f
.ends

.subckt PM_DFFLQNx1_ASAP7_75t_R%QN VSS 19 13 25 2 7 9 1 8
c1 1 VSS 0.00833483f
c2 2 VSS 0.00842221f
c3 7 VSS 0.00369824f
c4 8 VSS 0.00370094f
c5 9 VSS 0.00310013f
c6 10 VSS 0.00626829f
c7 11 VSS 0.00582839f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0115 $Y=0.2025 $X2=1.0240 $Y2=0.2025
r2 25 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0090 $Y=0.2025 $X2=1.0115 $Y2=0.2025
r3 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0260 $Y=0.2025
+ $X2=1.0260 $Y2=0.2340
r4 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.2340 $X2=1.0395 $Y2=0.2340
r5 11 20 1.09329 $w=1.76154e-08 $l=9.8e-09 $layer=M1 $thickness=3.6e-08
+ $X=1.0530 $Y=0.2340 $X2=1.0530 $Y2=0.2242
r6 11 23 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0530 $Y=0.2340 $X2=1.0395 $Y2=0.2340
r7 19 20 0.291487 $w=1.3e-08 $l=1.2e-09 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.2230 $X2=1.0530 $Y2=0.2242
r8 19 18 6.58761 $w=1.3e-08 $l=2.83e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.2230 $X2=1.0530 $Y2=0.1947
r9 17 18 15.4488 $w=1.3e-08 $l=6.62e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1285 $X2=1.0530 $Y2=0.1947
r10 9 16 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0530 $Y=0.0675 $X2=1.0530 $Y2=0.0360
r11 9 17 14.2246 $w=1.3e-08 $l=6.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.0675 $X2=1.0530 $Y2=0.1285
r12 15 16 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0395 $Y=0.0360 $X2=1.0530 $Y2=0.0360
r13 14 15 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.0360 $X2=1.0395 $Y2=0.0360
r14 10 14 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.0145
+ $Y=0.0360 $X2=1.0260 $Y2=0.0360
r15 1 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0260 $Y=0.0675
+ $X2=1.0260 $Y2=0.0360
r16 7 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.0115 $Y=0.0675 $X2=1.0240 $Y2=0.0675
r17 13 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.0090 $Y=0.0675 $X2=1.0115 $Y2=0.0675
.ends

.subckt PM_DFFLQNx1_ASAP7_75t_R%D VSS 9 3 4 1 6 5
c1 1 VSS 0.00677449f
c2 3 VSS 0.0834063f
c3 4 VSS 0.00583682f
c4 5 VSS 0.00681311f
c5 6 VSS 0.00761167f
r1 6 13 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.2340 $X2=0.2970 $Y2=0.2140
r2 5 8 5.17411 $w=1.46514e-08 $l=2.72e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0360 $X2=0.2970 $Y2=0.0632
r3 12 13 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1735 $X2=0.2970 $Y2=0.2140
r4 11 12 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1735
r5 9 10 2.85657 $w=1.3e-08 $l=1.22e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0820 $X2=0.2970 $Y2=0.0942
r6 9 8 4.37231 $w=1.3e-08 $l=1.88e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0820 $X2=0.2970 $Y2=0.0632
r7 4 10 5.07188 $w=1.3e-08 $l=2.18e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1160 $X2=0.2970 $Y2=0.0942
r8 4 11 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1160 $X2=0.2970 $Y2=0.1350
r9 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r10 1 11 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_DFFLQNx1_ASAP7_75t_R%CLK VSS 11 3 8 5 1 6 7 4
c1 1 VSS 0.00261925f
c2 3 VSS 0.0598036f
c3 4 VSS 0.00105358f
c4 5 VSS 0.00414449f
c5 6 VSS 0.00373881f
c6 7 VSS 0.00235168f
c7 8 VSS 0.00198947f
r1 6 17 3.22357 $w=2.26279e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.2125 $X2=0.1080 $Y2=0.1820
r2 5 15 3.22357 $w=2.26279e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0575 $X2=0.1080 $Y2=0.0880
r3 16 17 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.1820 $X2=0.1080 $Y2=0.1820
r4 8 13 2.6406 $w=2.38947e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1820 $X2=0.0810 $Y2=0.1540
r5 8 16 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1820 $X2=0.0945 $Y2=0.1820
r6 14 15 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.0880 $X2=0.1080 $Y2=0.0880
r7 7 10 1.76614 $w=2.65738e-08 $l=2.42e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0880 $X2=0.0810 $Y2=0.1122
r8 7 14 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0880 $X2=0.0945 $Y2=0.0880
r9 11 12 0.874462 $w=1.3e-08 $l=3.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1227
r10 11 10 1.57403 $w=1.3e-08 $l=6.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1122
r11 4 12 2.85657 $w=1.3e-08 $l=1.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1227
r12 4 13 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1540
r13 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r14 1 4 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_DFFLQNx1_ASAP7_75t_R%NET0109 VSS 2 4 1
c1 1 VSS 0.000984984f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0405 $X2=0.4905 $Y2=0.0405
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0405 $X2=0.4735 $Y2=0.0405
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4735 $Y=0.0405 $X2=0.4905 $Y2=0.0405
.ends

.subckt PM_DFFLQNx1_ASAP7_75t_R%NET06 VSS 2 4 1
c1 1 VSS 0.000973644f
r1 4 3 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3365 $Y2=0.2025
r2 2 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3195 $Y2=0.2025
r3 1 3 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3195 $Y=0.2025 $X2=0.3365 $Y2=0.2025
.ends

.subckt PM_DFFLQNx1_ASAP7_75t_R%NET0108 VSS 2 4 1
c1 1 VSS 0.000948527f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.2295 $X2=0.7605 $Y2=0.2295
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.2295 $X2=0.7435 $Y2=0.2295
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7435 $Y=0.2295 $X2=0.7605 $Y2=0.2295
.ends

.subckt PM_DFFLQNx1_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.00418102f
.ends

.subckt PM_DFFLQNx1_ASAP7_75t_R%NET0110 VSS 7 12 5 1 4
c1 1 VSS 0.00727636f
c2 4 VSS 0.00188706f
c3 5 VSS 0.00233436f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4880 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r3 9 5 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.4605
+ $Y=0.2295 $X2=0.4860 $Y2=0.2295
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.4455
+ $Y=0.2295 $X2=0.4605 $Y2=0.2295
r5 1 8 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4320
+ $Y=0.2295 $X2=0.4455 $Y2=0.2295
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2295 $X2=0.4300 $Y2=0.2295
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2295 $X2=0.4175 $Y2=0.2295
.ends

.subckt PM_DFFLQNx1_ASAP7_75t_R%NET020 VSS 7 10 5 4 1
c1 1 VSS 0.00972677f
c2 4 VSS 0.0031693f
c3 5 VSS 0.00186035f
r1 10 9 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r2 8 9 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r3 5 8 0.123457 $w=8.1e-08 $l=1e-08 $layer=N_src_drn $thickness=1e-09 $X=0.3780
+ $Y=0.0675 $X2=0.3880 $Y2=0.0675
r4 4 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3220 $Y2=0.0675
r5 7 4 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r6 1 5 1e-05
.ends

.subckt PM_DFFLQNx1_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.00417253f
.ends

.subckt PM_DFFLQNx1_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.00478249f
.ends

.subckt PM_DFFLQNx1_ASAP7_75t_R%NET0107 VSS 7 12 1 4 5
c1 1 VSS 0.00746711f
c2 4 VSS 0.00187637f
c3 5 VSS 0.00237802f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.0405 $X2=0.7705 $Y2=0.0405
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7580 $Y=0.0405 $X2=0.7705 $Y2=0.0405
r3 9 5 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.7425
+ $Y=0.0405 $X2=0.7560 $Y2=0.0405
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.7275
+ $Y=0.0405 $X2=0.7425 $Y2=0.0405
r5 1 8 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.7020
+ $Y=0.0405 $X2=0.7275 $Y2=0.0405
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.0405 $X2=0.7000 $Y2=0.0405
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.0405 $X2=0.6875 $Y2=0.0405
.ends

.subckt PM_DFFLQNx1_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.00470275f
.ends

.subckt PM_DFFLQNx1_ASAP7_75t_R%MH VSS 9 47 51 57 61 10 20 3 16 1 17 4 12 14 18
+ 15 19
c1 1 VSS 0.000275616f
c2 3 VSS 0.00624255f
c3 4 VSS 0.0054074f
c4 9 VSS 0.0363945f
c5 10 VSS 0.00226979f
c6 11 VSS 8.9782e-20
c7 12 VSS 0.00277968f
c8 13 VSS 6.86547e-20
c9 14 VSS 0.00851996f
c10 15 VSS 0.00125646f
c11 16 VSS 0.000667601f
c12 17 VSS 0.000550326f
c13 18 VSS 0.00649513f
c14 19 VSS 1.21068e-20
c15 20 VSS 0.00228255f
r1 61 60 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r2 59 60 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r3 3 59 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3760 $Y=0.2295 $X2=0.3880 $Y2=0.2295
r4 13 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2295 $X2=0.3760 $Y2=0.2295
r5 55 56 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r6 57 55 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.1890 $X2=0.3635 $Y2=0.1890
r7 12 56 0.185185 $w=5.4e-08 $l=1e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r8 12 3 0.518519 $w=3.9e-08 $l=4.05494e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.1890 $X2=0.3760 $Y2=0.2295
r9 3 44 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2295
+ $X2=0.3780 $Y2=0.2340
r10 51 50 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r11 49 50 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4420 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r12 4 49 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4300 $Y=0.0405 $X2=0.4420 $Y2=0.0405
r13 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0405 $X2=0.4300 $Y2=0.0405
r14 10 4 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0810 $X2=0.4300 $Y2=0.0810
r15 47 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0810 $X2=0.4175 $Y2=0.0810
r16 44 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r17 42 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r18 41 42 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4160
+ $Y=0.2340 $X2=0.4050 $Y2=0.2340
r19 14 20 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4340
+ $Y=0.2340 $X2=0.4590 $Y2=0.2340
r20 14 41 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4340
+ $Y=0.2340 $X2=0.4160 $Y2=0.2340
r21 4 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0405
+ $X2=0.4320 $Y2=0.0360
r22 20 34 3.01468 $w=1.741e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4590 $Y2=0.2140
r23 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4455 $Y2=0.0360
r24 18 31 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4590 $Y2=0.0630
r25 18 37 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4455 $Y2=0.0360
r26 33 34 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1850 $X2=0.4590 $Y2=0.2140
r27 32 33 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1660 $X2=0.4590 $Y2=0.1850
r28 16 19 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1525 $X2=0.4590 $Y2=0.1310
r29 16 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1525 $X2=0.4590 $Y2=0.1660
r30 30 31 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0900 $X2=0.4590 $Y2=0.0630
r31 29 30 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1025 $X2=0.4590 $Y2=0.0900
r32 15 19 2.78392 $w=1.56471e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1140 $X2=0.4590 $Y2=0.1310
r33 15 29 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1140 $X2=0.4590 $Y2=0.1025
r34 19 27 4.18306 $w=1.49565e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1310 $X2=0.4820 $Y2=0.1310
r35 26 27 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5000
+ $Y=0.1310 $X2=0.4820 $Y2=0.1310
r36 25 26 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1310 $X2=0.5000 $Y2=0.1310
r37 17 24 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1310 $X2=0.5670 $Y2=0.1310
r38 17 25 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1310 $X2=0.5130 $Y2=0.1310
r39 23 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1330
+ $X2=0.5670 $Y2=0.1310
r40 1 22 1.47681 $w=1.53e-08 $l=9e-09 $layer=LIG $thickness=4.8e-08 $X=0.5670
+ $Y=0.1215 $X2=0.5670 $Y2=0.1305
r41 22 23 5.31651 $w=1.53e-08 $l=2.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.5670 $Y=0.1305 $X2=0.5670 $Y2=0.1330
r42 9 22 0.314665 $w=2.27e-07 $l=4.5e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5670 $Y=0.1350 $X2=0.5670 $Y2=0.1305
r43 3 12 1e-05
.ends

.subckt PM_DFFLQNx1_ASAP7_75t_R%SS VSS 9 31 40 12 10 11 4 15 3 14 1 16 13 17
c1 1 VSS 0.00107388f
c2 3 VSS 0.00625652f
c3 4 VSS 0.00661555f
c4 9 VSS 0.0384305f
c5 10 VSS 0.00323747f
c6 11 VSS 0.00321889f
c7 12 VSS 0.00184572f
c8 13 VSS 0.0135797f
c9 14 VSS 0.0090072f
c10 15 VSS 0.00619013f
c11 16 VSS 0.00323823f
c12 17 VSS 0.00312873f
c13 18 VSS 0.00316228f
r1 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.2295 $X2=0.8620 $Y2=0.2295
r2 40 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.2295 $X2=0.8495 $Y2=0.2295
r3 4 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.2295
+ $X2=0.8640 $Y2=0.2340
r4 37 38 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.2340 $X2=0.8865 $Y2=0.2340
r5 14 18 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9180 $Y=0.2340 $X2=0.9450 $Y2=0.2340
r6 14 38 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.2340 $X2=0.8865 $Y2=0.2340
r7 18 35 6.74572 $w=1.545e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.2340 $X2=0.9450 $Y2=0.1980
r8 34 35 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1690 $X2=0.9450 $Y2=0.1980
r9 33 34 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1420 $X2=0.9450 $Y2=0.1690
r10 32 33 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1035 $X2=0.9450 $Y2=0.1420
r11 15 17 5.69636 $w=1.58e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.0675 $X2=0.9450 $Y2=0.0360
r12 15 32 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.0675 $X2=0.9450 $Y2=0.1035
r13 10 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.0405 $X2=0.8620 $Y2=0.0405
r14 31 10 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.0405 $X2=0.8495 $Y2=0.0405
r15 17 29 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.0360 $X2=0.9180 $Y2=0.0360
r16 3 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.0405
+ $X2=0.8640 $Y2=0.0360
r17 28 29 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.0360 $X2=0.9180 $Y2=0.0360
r18 27 28 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.0360 $X2=0.8910 $Y2=0.0360
r19 26 27 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.0360 $X2=0.8640 $Y2=0.0360
r20 13 16 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.0360 $X2=0.7830 $Y2=0.0360
r21 13 26 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0360 $X2=0.8370 $Y2=0.0360
r22 12 23 8.04505 $w=1.3e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.0705 $X2=0.7830 $Y2=0.1050
r23 12 16 6.39593 $w=1.55565e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7830 $Y=0.0705 $X2=0.7830 $Y2=0.0360
r24 1 20 2.36633 $w=2.3e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.7830
+ $Y=0.1055 $X2=0.7830 $Y2=0.1055
r25 1 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7830 $Y=0.1055
+ $X2=0.7830 $Y2=0.1050
r26 9 20 0.314665 $w=2.27e-07 $l=2.95e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.7830 $Y=0.1350 $X2=0.7830 $Y2=0.1055
.ends

.subckt PM_DFFLQNx1_ASAP7_75t_R%NET029 VSS 10 39 42 47 49 3 11 12 13 15 1 17 4
+ 18 14 16
c1 1 VSS 0.00219641f
c2 3 VSS 0.0053726f
c3 4 VSS 0.00934749f
c4 10 VSS 0.0374961f
c5 11 VSS 0.00286263f
c6 12 VSS 0.00269422f
c7 13 VSS 0.00225726f
c8 14 VSS 0.00186827f
c9 15 VSS 0.00403543f
c10 16 VSS 0.0029904f
c11 17 VSS 0.0010423f
c12 18 VSS 0.000415791f
c13 19 VSS 0.00295194f
r1 49 48 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.2295 $X2=0.6625 $Y2=0.2295
r2 13 48 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6500 $Y=0.2295 $X2=0.6625 $Y2=0.2295
r3 12 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2295 $X2=0.5920 $Y2=0.2295
r4 47 12 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.2295 $X2=0.5795 $Y2=0.2295
r5 44 13 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6210 $Y=0.2295 $X2=0.6480 $Y2=0.2295
r6 4 44 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08 $X=0.5940
+ $Y=0.2295 $X2=0.6210 $Y2=0.2295
r7 4 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2295
+ $X2=0.5965 $Y2=0.2340
r8 15 19 4.06404 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5965 $Y=0.2340 $X2=0.6210 $Y2=0.2340
r9 42 41 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.0405 $X2=0.6085 $Y2=0.0405
r10 40 41 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6040 $Y=0.0405 $X2=0.6085 $Y2=0.0405
r11 3 40 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5920 $Y=0.0405 $X2=0.6040 $Y2=0.0405
r12 11 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.0405 $X2=0.5920 $Y2=0.0405
r13 39 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0405 $X2=0.5795 $Y2=0.0405
r14 19 35 3.01468 $w=1.741e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.2340 $X2=0.6210 $Y2=0.2140
r15 3 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0405
+ $X2=0.5940 $Y2=0.0540
r16 34 35 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1850 $X2=0.6210 $Y2=0.2140
r17 33 34 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1660 $X2=0.6210 $Y2=0.1850
r18 32 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1525 $X2=0.6210 $Y2=0.1660
r19 31 32 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1310 $X2=0.6210 $Y2=0.1525
r20 17 28 3.60008 $w=1.51951e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.1105 $X2=0.6210 $Y2=0.0900
r21 17 31 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1105 $X2=0.6210 $Y2=0.1310
r22 16 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0540 $X2=0.5940 $Y2=0.0720
r23 27 28 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6075 $Y=0.0900 $X2=0.6210 $Y2=0.0900
r24 18 26 1.38478 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5940 $Y=0.0900 $X2=0.5830 $Y2=0.0900
r25 18 27 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5940 $Y=0.0900 $X2=0.6075 $Y2=0.0900
r26 18 29 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0900 $X2=0.5940 $Y2=0.0720
r27 25 26 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5515
+ $Y=0.0900 $X2=0.5830 $Y2=0.0900
r28 24 25 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0900 $X2=0.5515 $Y2=0.0900
r29 14 24 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5000
+ $Y=0.0900 $X2=0.5130 $Y2=0.0900
r30 1 21 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.5130
+ $Y=0.0900 $X2=0.5130 $Y2=0.0900
r31 1 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.0900
+ $X2=0.5130 $Y2=0.0900
r32 10 21 0.314665 $w=2.27e-07 $l=4.5e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5130 $Y2=0.0900
.ends

.subckt PM_DFFLQNx1_ASAP7_75t_R%CLKB VSS 11 12 57 59 17 6 5 16 15 13 21 22 14
+ 19 18 2 1 20
c1 1 VSS 4.23362e-20
c2 2 VSS 0.000131726f
c3 5 VSS 0.00727958f
c4 6 VSS 0.00729143f
c5 11 VSS 0.00437566f
c6 12 VSS 0.0045835f
c7 13 VSS 0.00648519f
c8 14 VSS 0.00649346f
c9 15 VSS 0.0102894f
c10 16 VSS 0.00855824f
c11 17 VSS 0.00622841f
c12 18 VSS 0.000546104f
c13 19 VSS 0.00156196f
c14 20 VSS 0.00361029f
c15 21 VSS 0.00300594f
c16 22 VSS 0.0168868f
r1 14 6 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1600 $Y2=0.2160
r2 59 14 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r3 13 5 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1600 $Y2=0.0540
r4 57 13 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r5 6 53 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r6 5 50 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r7 53 54 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1845 $Y2=0.2340
r8 16 21 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.2340 $X2=0.2430 $Y2=0.2340
r9 16 54 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.1845 $Y2=0.2340
r10 50 51 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1845 $Y2=0.0360
r11 15 20 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.0360 $X2=0.2430 $Y2=0.0360
r12 15 51 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.1845 $Y2=0.0360
r13 2 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6750 $Y=0.1350
+ $X2=0.6750 $Y2=0.1440
r14 12 2 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6750
+ $Y=0.1350 $X2=0.6750 $Y2=0.1350
r15 21 44 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.2340 $X2=0.2430 $Y2=0.2125
r16 20 41 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0360 $X2=0.2430 $Y2=0.0575
r17 19 45 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1125 $X2=0.6750 $Y2=0.1440
r18 43 44 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1990 $X2=0.2430 $Y2=0.2125
r19 42 43 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1890 $X2=0.2430 $Y2=0.1990
r20 40 41 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0880 $X2=0.2430 $Y2=0.0575
r21 39 40 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1160 $X2=0.2430 $Y2=0.0880
r22 38 42 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1710 $X2=0.2430 $Y2=0.1890
r23 37 38 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1530 $X2=0.2430 $Y2=0.1710
r24 17 37 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1530
r25 17 39 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1160
r26 35 45 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.6750 $Y=0.1530
+ $X2=0.6750 $Y2=0.1440
r27 34 35 18.3054 $w=1.3e-08 $l=7.85e-08 $layer=M2 $thickness=3.6e-08 $X=0.5965
+ $Y=0.1530 $X2=0.6750 $Y2=0.1530
r28 33 34 29.3819 $w=1.3e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.4705
+ $Y=0.1530 $X2=0.5965 $Y2=0.1530
r29 32 33 15.2739 $w=1.3e-08 $l=6.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1530 $X2=0.4705 $Y2=0.1530
r30 31 32 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1530 $X2=0.4050 $Y2=0.1530
r31 30 31 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1530 $X2=0.3240 $Y2=0.1530
r32 30 37 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.2430 $Y=0.1530
+ $X2=0.2430 $Y2=0.1530
r33 22 30 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.2315
+ $Y=0.1530 $X2=0.2430 $Y2=0.1530
r34 28 32 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4050 $Y=0.1440
+ $X2=0.4050 $Y2=0.1530
r35 18 28 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1160 $X2=0.4050 $Y2=0.1440
r36 11 1 5.63117 $w=1.26721e-07 $l=2e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4050 $Y2=0.1330
r37 1 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1330
+ $X2=0.4050 $Y2=0.1440
.ends

.subckt PM_DFFLQNx1_ASAP7_75t_R%SH VSS 11 12 59 62 65 68 14 23 25 13 6 18 16 17
+ 5 15 22 27 26 20 2 21 1 24 19 28
c1 1 VSS 0.000652967f
c2 2 VSS 0.00409702f
c3 5 VSS 0.00475822f
c4 6 VSS 0.00536486f
c5 11 VSS 0.0374658f
c6 12 VSS 0.0802607f
c7 13 VSS 0.0038063f
c8 14 VSS 0.00400055f
c9 15 VSS 0.00784986f
c10 16 VSS 0.00157811f
c11 17 VSS 0.00166999f
c12 18 VSS 0.00223064f
c13 19 VSS 0.000629172f
c14 20 VSS 0.000495232f
c15 21 VSS 0.00101611f
c16 22 VSS 0.00274731f
c17 23 VSS 0.00595729f
c18 24 VSS 0.00228357f
c19 25 VSS 0.000113837f
c20 26 VSS 0.000362455f
c21 27 VSS 0.000320625f
c22 28 VSS 0.00748195f
r1 68 67 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r2 5 67 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6500 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r3 64 5 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6380 $Y=0.0405 $X2=0.6500 $Y2=0.0405
r4 13 64 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0405 $X2=0.6380 $Y2=0.0405
r5 65 13 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.0405 $X2=0.6335 $Y2=0.0405
r6 62 61 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r7 60 61 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7120 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r8 6 60 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7000 $Y=0.2295 $X2=0.7120 $Y2=0.2295
r9 14 6 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.2295 $X2=0.7000 $Y2=0.2295
r10 59 14 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.2295 $X2=0.6875 $Y2=0.2295
r11 5 54 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.0405
+ $X2=0.6480 $Y2=0.0360
r12 2 49 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.9990 $Y=0.1350
+ $X2=0.9990 $Y2=0.1440
r13 12 2 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.9990
+ $Y=0.1350 $X2=0.9990 $Y2=0.1350
r14 6 47 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7020 $Y=0.2295
+ $X2=0.7020 $Y2=0.2340
r15 54 55 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6480
+ $Y=0.0360 $X2=0.6615 $Y2=0.0360
r16 52 55 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0360 $X2=0.6615 $Y2=0.0360
r17 51 52 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6860
+ $Y=0.0360 $X2=0.6750 $Y2=0.0360
r18 15 24 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.7040
+ $Y=0.0360 $X2=0.7290 $Y2=0.0360
r19 15 51 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7040
+ $Y=0.0360 $X2=0.6860 $Y2=0.0360
r20 22 49 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.9990
+ $Y=0.1080 $X2=0.9990 $Y2=0.1440
r21 47 48 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.2340 $X2=0.7155 $Y2=0.2340
r22 23 48 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.2340 $X2=0.7155 $Y2=0.2340
r23 24 40 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.0360 $X2=0.7290 $Y2=0.0630
r24 44 49 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.9990 $Y=0.1530
+ $X2=0.9990 $Y2=0.1440
r25 43 44 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1530 $X2=0.9990 $Y2=0.1530
r26 42 43 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1530 $X2=0.9450 $Y2=0.1530
r27 28 42 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.8795
+ $Y=0.1530 $X2=0.8910 $Y2=0.1530
r28 41 42 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.8910 $Y=0.1485 $X2=0.8910
+ $Y2=0.1530
r29 21 41 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1305 $X2=0.8910 $Y2=0.1485
r30 17 36 6.50021 $w=1.33448e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1980 $X2=0.7290 $Y2=0.1690
r31 17 23 7.21452 $w=1.425e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1980 $X2=0.7290 $Y2=0.2340
r32 39 40 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.0900 $X2=0.7290 $Y2=0.0630
r33 38 39 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1090 $X2=0.7290 $Y2=0.0900
r34 16 25 4.67854 $w=1.44583e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1360 $X2=0.7290 $Y2=0.1600
r35 16 38 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1360 $X2=0.7290 $Y2=0.1090
r36 27 37 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1575 $X2=0.8910 $Y2=0.1665
r37 27 41 1.50855 $w=1.55e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1575 $X2=0.8910 $Y2=0.1485
r38 27 42 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.8910 $Y=0.1575 $X2=0.8910
+ $Y2=0.1530
r39 25 36 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1600 $X2=0.7290 $Y2=0.1690
r40 35 37 4.19024 $w=1.156e-08 $l=2.54018e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8660 $Y=0.1620 $X2=0.8910 $Y2=0.1665
r41 20 26 1.38478 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8480 $Y=0.1620 $X2=0.8370 $Y2=0.1620
r42 20 35 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8480
+ $Y=0.1620 $X2=0.8660 $Y2=0.1620
r43 34 36 4.4015 $w=1.35e-08 $l=2.78927e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7560 $Y=0.1620 $X2=0.7290 $Y2=0.1690
r44 33 34 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1620 $X2=0.7560 $Y2=0.1620
r45 18 26 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.1620 $X2=0.8370 $Y2=0.1620
r46 18 33 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.1620 $X2=0.7830 $Y2=0.1620
r47 26 32 4.88263 $w=1.47308e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8370 $Y=0.1620 $X2=0.8370 $Y2=0.1360
r48 19 32 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1180 $X2=0.8370 $Y2=0.1360
r49 11 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.8370
+ $Y=0.1350 $X2=0.8370 $Y2=0.1350
r50 1 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8370 $Y=0.1350
+ $X2=0.8370 $Y2=0.1360
.ends

.subckt PM_DFFLQNx1_ASAP7_75t_R%CLKN VSS 16 17 18 19 20 99 101 28 35 32 9 34 8
+ 21 22 26 25 1 27 36 23 29 2 5 30 3 10 31 33 24
c1 1 VSS 0.00148342f
c2 2 VSS 0.000298569f
c3 3 VSS 7.25042e-20
c4 4 VSS 1e-36
c5 5 VSS 0.000412174f
c6 8 VSS 0.00771313f
c7 9 VSS 0.00771726f
c8 10 VSS 0.00355108f
c9 16 VSS 0.0590851f
c10 17 VSS 0.00560537f
c11 18 VSS 0.0051156f
c12 19 VSS 0.00437881f
c13 20 VSS 0.00517314f
c14 21 VSS 0.00655762f
c15 22 VSS 0.00650818f
c16 23 VSS 0.00804272f
c17 24 VSS 0.00180719f
c18 25 VSS 0.00454152f
c19 26 VSS 0.00375638f
c20 27 VSS 0.000658378f
c21 28 VSS 0.000261282f
c22 29 VSS 0.000826989f
c23 30 VSS 0.00146331f
c24 31 VSS 0.00383175f
c25 32 VSS 0.00190563f
c26 33 VSS 0.00393268f
c27 34 VSS 0.00084138f
c28 35 VSS 0.000477266f
c29 36 VSS 0.0229229f
r1 101 100 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r2 22 100 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r3 99 98 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r4 21 98 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r5 9 96 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0550 $Y2=0.2340
r6 8 93 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0550 $Y2=0.0360
r7 95 96 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.2340 $X2=0.0550 $Y2=0.2340
r8 26 95 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0460 $Y2=0.2340
r9 26 33 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0180 $Y2=0.2340
r10 92 93 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.0360 $X2=0.0550 $Y2=0.0360
r11 25 92 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0460 $Y2=0.0360
r12 25 31 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0180 $Y2=0.0360
r13 5 91 2.78395 $w=2.4e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08 $X=0.7290
+ $Y=0.1780 $X2=0.7250 $Y2=0.1780
r14 20 5 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.7290 $Y=0.1350 $X2=0.7290 $Y2=0.1780
r15 4 84 10.3807 $w=2.30357e-08 $l=0 $layer=LISD $thickness=3.675e-08 $X=0.6210
+ $Y=0.1780 $X2=0.6210 $Y2=0.1780
r16 19 4 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.6210 $Y=0.1350 $X2=0.6210 $Y2=0.1780
r17 3 77 2.78395 $w=2.4e-08 $l=5e-09 $layer=LIG $thickness=4.8e-08 $X=0.4590
+ $Y=0.1780 $X2=0.4640 $Y2=0.1780
r18 18 3 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4590 $Y2=0.1780
r19 33 72 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.2340 $X2=0.0180 $Y2=0.2125
r20 31 71 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.0360 $X2=0.0180 $Y2=0.0575
r21 90 91 4.8113 $w=2.22e-08 $l=1.5e-09 $layer=LISD $thickness=2.7e-08
+ $X=0.7235 $Y=0.1780 $X2=0.7250 $Y2=0.1780
r22 89 90 10.8887 $w=2.22e-08 $l=2.15e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7020 $Y=0.1780 $X2=0.7235 $Y2=0.1780
r23 88 89 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6885 $Y=0.1780 $X2=0.7020 $Y2=0.1780
r24 87 88 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6750 $Y=0.1780 $X2=0.6885 $Y2=0.1780
r25 86 87 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6615 $Y=0.1780 $X2=0.6750 $Y2=0.1780
r26 85 86 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6480 $Y=0.1780 $X2=0.6615 $Y2=0.1780
r27 84 85 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6210 $Y=0.1780 $X2=0.6480 $Y2=0.1780
r28 83 84 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5940 $Y=0.1780 $X2=0.6210 $Y2=0.1780
r29 82 83 7.09034 $w=2.22e-08 $l=1.4e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5800 $Y=0.1780 $X2=0.5940 $Y2=0.1780
r30 81 82 6.58388 $w=2.22e-08 $l=1.3e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5670 $Y=0.1780 $X2=0.5800 $Y2=0.1780
r31 80 81 6.58388 $w=2.22e-08 $l=1.3e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5540 $Y=0.1780 $X2=0.5670 $Y2=0.1780
r32 79 80 7.09034 $w=2.22e-08 $l=1.4e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5400 $Y=0.1780 $X2=0.5540 $Y2=0.1780
r33 78 79 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5265 $Y=0.1780 $X2=0.5400 $Y2=0.1780
r34 76 77 10.3823 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4775 $Y=0.1780 $X2=0.4640 $Y2=0.1780
r35 75 76 11.142 $w=2.22e-08 $l=2.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4995 $Y=0.1780 $X2=0.4775 $Y2=0.1780
r36 74 78 1.51936 $w=2.22e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.5235
+ $Y=0.1780 $X2=0.5265 $Y2=0.1780
r37 73 74 5.31775 $w=2.22e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5130 $Y=0.1780 $X2=0.5235 $Y2=0.1780
r38 10 73 5.31775 $w=2.22e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5025 $Y=0.1780 $X2=0.5130 $Y2=0.1780
r39 10 75 1.51936 $w=2.22e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.5025
+ $Y=0.1780 $X2=0.4995 $Y2=0.1780
r40 2 65 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
r41 17 2 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r42 24 32 0.998523 $w=1.74118e-08 $l=1.01119e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1990 $X2=0.0165 $Y2=0.1890
r43 24 72 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1990 $X2=0.0180 $Y2=0.2125
r44 70 71 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0880 $X2=0.0180 $Y2=0.0575
r45 69 70 10.9599 $w=1.3e-08 $l=4.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1350 $X2=0.0180 $Y2=0.0880
r46 23 32 2.63085 $w=1.54194e-08 $l=1.7066e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1720 $X2=0.0165 $Y2=0.1890
r47 23 69 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1720 $X2=0.0180 $Y2=0.1350
r48 67 73 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5130 $Y=0.1845
+ $X2=0.5130 $Y2=0.1780
r49 30 67 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1680 $X2=0.5130 $Y2=0.1845
r50 65 66 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1555
r51 29 63 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1735 $X2=0.3510 $Y2=0.1890
r52 29 66 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1735 $X2=0.3510 $Y2=0.1555
r53 60 61 1.90199 $w=1.38333e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.0255 $Y=0.1890 $X2=0.0345 $Y2=0.1890
r54 32 60 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0165
+ $Y=0.1890 $X2=0.0255 $Y2=0.1890
r55 58 67 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.5130 $Y=0.1890
+ $X2=0.5130 $Y2=0.1845
r56 57 58 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.4320
+ $Y=0.1890 $X2=0.5130 $Y2=0.1890
r57 56 57 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1890 $X2=0.4320 $Y2=0.1890
r58 56 63 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.3510 $Y=0.1890
+ $X2=0.3510 $Y2=0.1890
r59 55 56 15.2739 $w=1.3e-08 $l=6.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.2855
+ $Y=0.1890 $X2=0.3510 $Y2=0.1890
r60 54 55 20.2875 $w=1.3e-08 $l=8.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.1985
+ $Y=0.1890 $X2=0.2855 $Y2=0.1890
r61 53 54 9.211 $w=1.3e-08 $l=3.95e-08 $layer=M2 $thickness=3.6e-08 $X=0.1590
+ $Y=0.1890 $X2=0.1985 $Y2=0.1890
r62 52 53 14.691 $w=1.3e-08 $l=6.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.0960
+ $Y=0.1890 $X2=0.1590 $Y2=0.1890
r63 51 52 14.691 $w=1.3e-08 $l=6.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.0330
+ $Y=0.1890 $X2=0.0960 $Y2=0.1890
r64 51 61 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.0330 $Y=0.1890
+ $X2=0.0345 $Y2=0.1890
r65 36 51 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.0215
+ $Y=0.1890 $X2=0.0330 $Y2=0.1890
r66 48 49 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1590
+ $Y=0.1890 $X2=0.1740 $Y2=0.1890
r67 48 53 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1590 $Y=0.1890
+ $X2=0.1590 $Y2=0.1890
r68 34 46 2.78392 $w=1.56471e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1890 $X2=0.1890 $Y2=0.1720
r69 34 49 2.31754 $w=1.6e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1890 $X2=0.1740 $Y2=0.1890
r70 28 35 2.78149 $w=1.76421e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1540 $X2=0.1890 $Y2=0.1350
r71 28 46 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1540 $X2=0.1890 $Y2=0.1720
r72 35 45 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1640 $Y2=0.1350
r73 44 45 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.1465
+ $Y=0.1350 $X2=0.1640 $Y2=0.1350
r74 43 44 0.46638 $w=1.3e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.1445
+ $Y=0.1350 $X2=0.1465 $Y2=0.1350
r75 42 43 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1445 $Y2=0.1350
r76 27 42 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1235
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r77 16 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r78 1 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
r79 9 22 1e-05
r80 8 21 1e-05
.ends


*
.SUBCKT DFFLQNx1_ASAP7_75t_R VSS VDD CLK D QN
*
* VSS VSS
* VDD VDD
* CLK CLK
* D D
* QN QN
*
*

MM20 N_MM20_d N_MM20_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM23 N_MM23_d N_MM22_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM10_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM6 N_MM6_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM12 N_MM12_d N_MM12_g N_MM12_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM17 N_MM17_d N_MM13_g N_MM17_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM16 N_MM16_d N_MM19_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM14 N_MM14_d N_MM14_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM24 N_MM24_d N_MM24_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM21 N_MM21_d N_MM20_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM22 N_MM22_d N_MM22_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM13 N_MM13_d N_MM13_g N_MM13_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM18 N_MM18_d N_MM18_g N_MM18_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM19 N_MM19_d N_MM19_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM15 N_MM15_d N_MM14_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM25 N_MM25_d N_MM24_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "DFFLQNx1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "DFFLQNx1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_DFFLQNx1_ASAP7_75t_R%noxref_29 VSS N_noxref_29_1
+ PM_DFFLQNx1_ASAP7_75t_R%noxref_29
cc_1 N_noxref_29_1 N_MM24_g 0.00148755f
cc_2 N_noxref_29_1 N_QN_8 0.0385769f
cc_3 N_noxref_29_1 N_noxref_28_1 0.00177063f
x_PM_DFFLQNx1_ASAP7_75t_R%noxref_28 VSS N_noxref_28_1
+ PM_DFFLQNx1_ASAP7_75t_R%noxref_28
cc_4 N_noxref_28_1 N_MM24_g 0.00148752f
cc_5 N_noxref_28_1 N_QN_7 0.0383585f
x_PM_DFFLQNx1_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_DFFLQNx1_ASAP7_75t_R%noxref_22
cc_6 N_noxref_22_1 N_MM3_g 0.00136567f
cc_7 N_noxref_22_1 N_CLKB_13 0.000803613f
cc_8 N_noxref_22_1 N_noxref_20_1 0.00770008f
cc_9 N_noxref_22_1 N_noxref_21_1 0.000471857f
x_PM_DFFLQNx1_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_DFFLQNx1_ASAP7_75t_R%noxref_23
cc_10 N_noxref_23_1 N_MM3_g 0.00137373f
cc_11 N_noxref_23_1 N_CLKB_14 0.000769423f
cc_12 N_noxref_23_1 N_noxref_20_1 0.000469294f
cc_13 N_noxref_23_1 N_noxref_21_1 0.00769869f
cc_14 N_noxref_23_1 N_noxref_22_1 0.00123383f
x_PM_DFFLQNx1_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_DFFLQNx1_ASAP7_75t_R%noxref_24
cc_15 N_noxref_24_1 N_SS_10 0.0170238f
cc_16 N_noxref_24_1 N_MM14_g 0.00611563f
x_PM_DFFLQNx1_ASAP7_75t_R%noxref_26 VSS N_noxref_26_1
+ PM_DFFLQNx1_ASAP7_75t_R%noxref_26
cc_17 N_noxref_26_1 N_SS_10 0.00063571f
cc_18 N_noxref_26_1 N_MM24_g 0.0016864f
cc_19 N_noxref_26_1 N_noxref_24_1 0.00776266f
cc_20 N_noxref_26_1 N_noxref_25_1 0.0004811f
x_PM_DFFLQNx1_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_DFFLQNx1_ASAP7_75t_R%noxref_25
cc_21 N_noxref_25_1 N_SS_11 0.0168754f
cc_22 N_noxref_25_1 N_SH_1 0.000168104f
cc_23 N_noxref_25_1 N_MM14_g 0.00601738f
cc_24 N_noxref_25_1 N_noxref_24_1 0.00153369f
x_PM_DFFLQNx1_ASAP7_75t_R%noxref_27 VSS N_noxref_27_1
+ PM_DFFLQNx1_ASAP7_75t_R%noxref_27
cc_25 N_noxref_27_1 N_SS_11 0.000625524f
cc_26 N_noxref_27_1 N_MM24_g 0.00170724f
cc_27 N_noxref_27_1 N_noxref_24_1 0.000482678f
cc_28 N_noxref_27_1 N_noxref_25_1 0.00776535f
cc_29 N_noxref_27_1 N_noxref_26_1 0.00124093f
x_PM_DFFLQNx1_ASAP7_75t_R%QN VSS QN N_MM24_d N_MM25_d N_QN_2 N_QN_7 N_QN_9
+ N_QN_1 N_QN_8 PM_DFFLQNx1_ASAP7_75t_R%QN
cc_30 N_QN_2 N_SS_17 0.000428924f
cc_31 N_QN_2 N_SS_15 0.00179586f
cc_32 N_QN_7 N_SH_22 0.00111416f
cc_33 N_QN_9 N_SH_28 0.000793765f
cc_34 N_QN_2 N_SH_2 0.000895953f
cc_35 N_QN_2 N_MM24_g 0.0011755f
cc_36 N_QN_1 N_MM24_g 0.0012462f
cc_37 N_QN_8 N_SH_2 0.00157238f
cc_38 N_QN_9 N_SH_22 0.00540121f
cc_39 N_QN_8 N_MM24_g 0.015456f
cc_40 N_QN_7 N_MM24_g 0.0543696f
x_PM_DFFLQNx1_ASAP7_75t_R%D VSS D N_MM3_g N_D_4 N_D_1 N_D_6 N_D_5
+ PM_DFFLQNx1_ASAP7_75t_R%D
cc_41 N_MM3_g N_CLKN_29 0.000914141f
cc_42 N_D_4 N_CLKN_36 0.000997257f
cc_43 N_D_1 N_CLKN_2 0.00239967f
cc_44 N_D_4 N_CLKN_29 0.00461054f
cc_45 N_MM3_g N_MM1_g 0.00527302f
x_PM_DFFLQNx1_ASAP7_75t_R%CLK VSS CLK N_MM20_g N_CLK_8 N_CLK_5 N_CLK_1 N_CLK_6
+ N_CLK_7 N_CLK_4 PM_DFFLQNx1_ASAP7_75t_R%CLK
x_PM_DFFLQNx1_ASAP7_75t_R%NET0109 VSS N_MM9_s N_MM8_d N_NET0109_1
+ PM_DFFLQNx1_ASAP7_75t_R%NET0109
cc_46 N_NET0109_1 N_MM9_g 0.00772304f
cc_47 N_NET0109_1 N_MM11_g 0.00772856f
x_PM_DFFLQNx1_ASAP7_75t_R%NET06 VSS N_MM3_d N_MM1_s N_NET06_1
+ PM_DFFLQNx1_ASAP7_75t_R%NET06
cc_48 N_NET06_1 N_MM1_g 0.0169405f
cc_49 N_NET06_1 N_MM3_g 0.0170094f
x_PM_DFFLQNx1_ASAP7_75t_R%NET0108 VSS N_MM18_s N_MM19_d N_NET0108_1
+ PM_DFFLQNx1_ASAP7_75t_R%NET0108
cc_50 N_NET0108_1 N_MM18_g 0.00773054f
cc_51 N_NET0108_1 N_MM19_g 0.00776247f
x_PM_DFFLQNx1_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_DFFLQNx1_ASAP7_75t_R%noxref_18
cc_52 N_noxref_18_1 N_MM20_g 0.00368833f
cc_53 N_noxref_18_1 N_CLKN_8 0.000543714f
cc_54 N_noxref_18_1 N_CLKN_9 4.21487e-20
cc_55 N_noxref_18_1 N_CLKN_31 5.87338e-20
cc_56 N_noxref_18_1 N_CLKN_23 0.000384924f
cc_57 N_noxref_18_1 N_CLKN_21 0.0276297f
x_PM_DFFLQNx1_ASAP7_75t_R%NET0110 VSS N_MM10_s N_MM11_d N_NET0110_5 N_NET0110_1
+ N_NET0110_4 PM_DFFLQNx1_ASAP7_75t_R%NET0110
cc_58 N_NET0110_5 N_CLKN_10 0.00146263f
cc_59 N_NET0110_1 N_CLKN_3 0.00052085f
cc_60 N_NET0110_1 N_MM9_g 0.00206401f
cc_61 N_NET0110_4 N_MM9_g 0.00714445f
cc_62 N_NET0110_5 N_MM9_g 0.0240626f
cc_63 N_NET0110_4 N_MM10_g 0.0150104f
cc_64 N_NET0110_5 N_MM11_g 0.0145937f
cc_65 N_NET0110_1 N_MH_16 0.000461869f
cc_66 N_NET0110_4 N_MH_3 0.000601242f
cc_67 N_NET0110_1 N_MH_20 0.00323624f
x_PM_DFFLQNx1_ASAP7_75t_R%NET020 VSS N_MM5_d N_MM4_s N_NET020_5 N_NET020_4
+ N_NET020_1 PM_DFFLQNx1_ASAP7_75t_R%NET020
cc_68 N_NET020_5 N_CLKN_29 0.000206755f
cc_69 N_NET020_5 N_CLKN_2 0.0020947f
cc_70 N_NET020_5 N_MM1_g 0.0733026f
cc_71 N_NET020_4 N_D_1 0.000671161f
cc_72 N_NET020_4 N_D_4 0.00076378f
cc_73 N_NET020_4 N_MM3_g 0.0361889f
cc_74 N_NET020_5 N_CLKB_18 0.000306104f
cc_75 N_NET020_5 N_CLKB_1 0.000757233f
cc_76 N_NET020_5 N_MM10_g 0.0346066f
cc_77 N_NET020_1 N_MH_4 0.00121047f
cc_78 N_NET020_1 N_MH_10 0.00348758f
x_PM_DFFLQNx1_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_DFFLQNx1_ASAP7_75t_R%noxref_19
cc_79 N_noxref_19_1 N_MM20_g 0.00367454f
cc_80 N_noxref_19_1 N_CLKN_8 4.38676e-20
cc_81 N_noxref_19_1 N_CLKN_33 5.38656e-20
cc_82 N_noxref_19_1 N_CLKN_24 8.26328e-20
cc_83 N_noxref_19_1 N_CLKN_32 8.8491e-20
cc_84 N_noxref_19_1 N_CLKN_23 0.000272497f
cc_85 N_noxref_19_1 N_CLKN_9 0.00050327f
cc_86 N_noxref_19_1 N_CLKN_22 0.0277397f
cc_87 N_noxref_19_1 N_noxref_18_1 0.00204446f
x_PM_DFFLQNx1_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_DFFLQNx1_ASAP7_75t_R%noxref_20
cc_88 N_noxref_20_1 N_CLKN_1 0.000129137f
cc_89 N_noxref_20_1 N_MM22_g 0.00352737f
cc_90 N_noxref_20_1 N_CLKB_5 0.000443316f
cc_91 N_noxref_20_1 N_CLKB_13 0.0271662f
x_PM_DFFLQNx1_ASAP7_75t_R%NET0107 VSS N_MM17_s N_MM16_d N_NET0107_1 N_NET0107_4
+ N_NET0107_5 PM_DFFLQNx1_ASAP7_75t_R%NET0107
cc_92 N_NET0107_1 N_MM18_g 0.000859473f
cc_93 N_NET0107_4 N_MM18_g 0.00695814f
cc_94 N_NET0107_5 N_MM18_g 0.0240007f
cc_95 N_NET0107_4 N_MM13_g 0.0153014f
cc_96 N_NET0107_1 N_MM19_g 0.000917747f
cc_97 N_NET0107_5 N_MM19_g 0.0155804f
cc_98 N_NET0107_1 N_SH_13 0.000516418f
cc_99 N_NET0107_1 N_SH_15 0.000461115f
cc_100 N_NET0107_1 N_SH_16 0.000600253f
cc_101 N_NET0107_4 N_SH_5 0.000661866f
cc_102 N_NET0107_1 N_SH_24 0.00237063f
x_PM_DFFLQNx1_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_DFFLQNx1_ASAP7_75t_R%noxref_21
cc_103 N_noxref_21_1 N_CLKN_1 0.000125863f
cc_104 N_noxref_21_1 N_MM22_g 0.00366742f
cc_105 N_noxref_21_1 N_CLKB_6 0.000435904f
cc_106 N_noxref_21_1 N_CLKB_14 0.0270926f
cc_107 N_noxref_21_1 N_noxref_20_1 0.00146986f
x_PM_DFFLQNx1_ASAP7_75t_R%MH VSS N_MM7_g N_MM4_d N_MM9_d N_MM1_d N_MM10_d
+ N_MH_10 N_MH_20 N_MH_3 N_MH_16 N_MH_1 N_MH_17 N_MH_4 N_MH_12 N_MH_14 N_MH_18
+ N_MH_15 N_MH_19 PM_DFFLQNx1_ASAP7_75t_R%MH
cc_108 N_MH_10 N_CLKN_30 0.000373765f
cc_109 N_MH_10 N_MM1_g 0.00040242f
cc_110 N_MH_10 N_CLKN_29 0.000392224f
cc_111 N_MH_20 N_CLKN_30 0.000254821f
cc_112 N_MH_3 N_CLKN_2 0.000280434f
cc_113 N_MH_16 N_CLKN_30 0.00268657f
cc_114 N_MH_1 N_CLKN_10 0.00208787f
cc_115 N_MH_17 N_CLKN_10 0.000621023f
cc_116 N_MH_4 N_MM9_g 0.000631784f
cc_117 N_MH_16 N_CLKN_3 0.000763461f
cc_118 N_MH_12 N_CLKN_2 0.000880682f
cc_119 N_MH_3 N_CLKN_29 0.00133137f
cc_120 N_MH_14 N_CLKN_29 0.00140466f
cc_121 N_MH_14 N_CLKN_36 0.00151046f
cc_122 N_MH_3 N_MM1_g 0.0017757f
cc_123 N_MH_17 N_CLKN_30 0.0036172f
cc_124 N_MM7_g N_CLKN_10 0.00459974f
cc_125 N_MH_12 N_MM1_g 0.0337007f
cc_126 N_MM7_g N_MM12_g 0.0127497f
cc_127 N_MH_10 N_MM9_g 0.0363082f
cc_128 N_MH_10 N_MM13_g 0.000161633f
cc_129 N_MH_10 N_CLKB_18 0.000266058f
cc_130 N_MH_14 N_CLKB_18 0.000329883f
cc_131 N_MH_18 N_CLKB_18 0.000380639f
cc_132 N_MH_12 N_MM10_g 0.016421f
cc_133 N_MH_3 N_CLKB_1 0.000736168f
cc_134 N_MH_4 N_MM10_g 0.00109525f
cc_135 N_MH_15 N_CLKB_18 0.00111823f
cc_136 N_MH_3 N_MM10_g 0.0011739f
cc_137 N_MH_17 N_CLKB_22 0.00124911f
cc_138 N_MH_16 N_CLKB_18 0.00135159f
cc_139 N_MH_12 N_CLKB_1 0.00182497f
cc_140 N_MH_16 N_CLKB_22 0.00230074f
cc_141 N_MH_19 N_CLKB_18 0.00273106f
cc_142 N_MH_10 N_MM10_g 0.0530757f
cc_143 N_MH_4 N_NET029_1 0.000401736f
cc_144 N_MH_17 N_NET029_18 0.000563962f
cc_145 N_MH_17 N_NET029_1 0.00083004f
cc_146 N_MH_1 N_NET029_14 0.000836245f
cc_147 N_MM7_g N_NET029_3 0.000974704f
cc_148 N_MH_17 N_NET029_17 0.00100361f
cc_149 N_MH_1 N_MM11_g 0.00106062f
cc_150 N_MM7_g N_NET029_1 0.00116078f
cc_151 N_MH_15 N_NET029_14 0.00123984f
cc_152 N_MM7_g N_NET029_12 0.00639534f
cc_153 N_MM7_g N_NET029_11 0.0064086f
cc_154 N_MH_17 N_NET029_14 0.00719398f
cc_155 N_MM7_g N_MM11_g 0.0293026f
x_PM_DFFLQNx1_ASAP7_75t_R%SS VSS N_MM19_g N_MM14_d N_MM15_d N_SS_12 N_SS_10
+ N_SS_11 N_SS_4 N_SS_15 N_SS_3 N_SS_14 N_SS_1 N_SS_16 N_SS_13 N_SS_17
+ PM_DFFLQNx1_ASAP7_75t_R%SS
cc_156 N_MM19_g N_CLKN_10 0.000218803f
cc_157 N_MM19_g N_CLKN_5 0.000537557f
cc_158 N_MM19_g N_MM18_g 0.013531f
x_PM_DFFLQNx1_ASAP7_75t_R%NET029 VSS N_MM11_g N_MM6_d N_MM12_d N_MM7_d N_MM13_d
+ N_NET029_3 N_NET029_11 N_NET029_12 N_NET029_13 N_NET029_15 N_NET029_1
+ N_NET029_17 N_NET029_4 N_NET029_18 N_NET029_14 N_NET029_16
+ PM_DFFLQNx1_ASAP7_75t_R%NET029
cc_159 N_NET029_3 N_CLKN_30 0.000491884f
cc_160 N_NET029_3 N_CLKN_10 0.000583014f
cc_161 N_NET029_3 N_CLKN_3 0.000123997f
cc_162 N_NET029_3 N_MM9_g 0.000162223f
cc_163 N_NET029_3 N_CLKN_36 0.000189583f
cc_164 N_NET029_11 N_MM12_g 0.00678159f
cc_165 N_NET029_12 N_MM12_g 0.00780029f
cc_166 N_NET029_13 N_MM12_g 0.00777313f
cc_167 N_NET029_15 N_CLKN_10 0.00037499f
cc_168 N_NET029_1 N_MM9_g 0.000568367f
cc_169 N_NET029_17 N_CLKN_10 0.00155422f
cc_170 N_NET029_4 N_MM12_g 0.00231951f
cc_171 N_NET029_4 N_CLKN_10 0.00634492f
cc_172 N_MM11_g N_MM9_g 0.0143808f
cc_173 N_NET029_3 N_MM12_g 0.0257229f
cc_174 N_NET029_13 N_MM10_g 0.000130173f
cc_175 N_NET029_13 N_CLKB_19 0.000373467f
cc_176 N_NET029_13 N_CLKB_22 0.000205442f
cc_177 N_NET029_13 N_CLKB_2 0.000228023f
cc_178 N_NET029_17 N_CLKB_19 0.00440577f
cc_179 N_NET029_17 N_CLKB_2 0.000385636f
cc_180 N_NET029_18 N_CLKB_19 0.00066483f
cc_181 N_NET029_14 N_CLKB_22 0.00268775f
cc_182 N_NET029_13 N_MM13_g 0.0153918f
x_PM_DFFLQNx1_ASAP7_75t_R%CLKB VSS N_MM10_g N_MM13_g N_MM23_d N_MM22_d
+ N_CLKB_17 N_CLKB_6 N_CLKB_5 N_CLKB_16 N_CLKB_15 N_CLKB_13 N_CLKB_21 N_CLKB_22
+ N_CLKB_14 N_CLKB_19 N_CLKB_18 N_CLKB_2 N_CLKB_1 N_CLKB_20
+ PM_DFFLQNx1_ASAP7_75t_R%CLKB
cc_183 N_CLKB_17 N_CLK_5 9.42407e-20
cc_184 N_CLKB_6 N_CLK_5 0.000321239f
cc_185 N_CLKB_5 N_CLK_5 0.000406233f
cc_186 N_CLKB_16 N_CLK_5 0.000213606f
cc_187 N_CLKB_16 N_CLK_6 0.000974336f
cc_188 N_CLKB_15 N_CLK_5 0.00219578f
cc_189 N_CLKB_13 N_CLKN_26 3.22363e-20
cc_190 N_CLKB_13 N_CLKN_23 6.25695e-20
cc_191 N_MM13_g N_CLKN_5 0.000222584f
cc_192 N_CLKB_21 N_CLKN_34 0.000231065f
cc_193 N_CLKB_6 N_CLKN_34 0.000271072f
cc_194 N_CLKB_22 N_CLKN_30 0.000665549f
cc_195 N_CLKB_6 N_CLKN_1 0.000308943f
cc_196 N_CLKB_14 N_MM22_g 0.0112471f
cc_197 N_CLKB_16 N_CLKN_34 0.00508495f
cc_198 N_CLKB_22 N_CLKN_29 0.000355479f
cc_199 N_CLKB_15 N_CLKN_35 0.000485317f
cc_200 N_MM10_g N_CLKN_3 0.000540881f
cc_201 N_CLKB_19 N_CLKN_10 0.000573169f
cc_202 N_CLKB_18 N_CLKN_36 0.000611247f
cc_203 N_CLKB_14 N_CLKN_1 0.000622622f
cc_204 N_CLKB_6 N_CLKN_27 0.000664076f
cc_205 N_CLKB_2 N_CLKN_10 0.00285577f
cc_206 N_CLKB_17 N_CLKN_36 0.000735061f
cc_207 N_CLKB_5 N_MM22_g 0.000758246f
cc_208 N_CLKB_1 N_CLKN_2 0.00227225f
cc_209 N_CLKB_17 N_CLKN_28 0.000987161f
cc_210 N_CLKB_6 N_MM22_g 0.00107449f
cc_211 N_MM10_g N_MM1_g 0.00163138f
cc_212 N_CLKB_18 N_CLKN_29 0.00310318f
cc_213 N_CLKB_17 N_CLKN_35 0.00376568f
cc_214 N_MM13_g N_CLKN_10 0.00430634f
cc_215 N_MM13_g N_MM12_g 0.00567097f
cc_216 N_MM10_g N_MM9_g 0.00910718f
cc_217 N_MM13_g N_MM18_g 0.0184479f
cc_218 N_CLKB_22 N_CLKN_36 0.0284489f
cc_219 N_CLKB_13 N_MM22_g 0.03884f
cc_220 N_CLKB_18 N_D_4 0.000146015f
cc_221 N_CLKB_21 N_D_6 0.000777105f
cc_222 N_CLKB_20 N_D_5 0.00096655f
cc_223 N_CLKB_22 N_D_4 0.00114922f
cc_224 N_CLKB_17 N_D_4 0.00840474f
x_PM_DFFLQNx1_ASAP7_75t_R%SH VSS N_MM14_g N_MM24_g N_MM13_s N_MM18_d N_MM12_s
+ N_MM17_d N_SH_14 N_SH_23 N_SH_25 N_SH_13 N_SH_6 N_SH_18 N_SH_16 N_SH_17
+ N_SH_5 N_SH_15 N_SH_22 N_SH_27 N_SH_26 N_SH_20 N_SH_2 N_SH_21 N_SH_1 N_SH_24
+ N_SH_19 N_SH_28 PM_DFFLQNx1_ASAP7_75t_R%SH
cc_225 N_SH_14 N_CLKN_36 9.89119e-20
cc_226 N_SH_23 N_CLKN_10 0.000170657f
cc_227 N_SH_25 N_CLKN_10 0.000204456f
cc_228 N_SH_13 N_MM12_g 0.00677846f
cc_229 N_SH_6 N_CLKN_10 0.000267105f
cc_230 N_SH_18 N_CLKN_5 0.000408984f
cc_231 N_SH_16 N_CLKN_10 0.000419671f
cc_232 N_SH_17 N_CLKN_10 0.000588129f
cc_233 N_SH_14 N_CLKN_5 0.000929177f
cc_234 N_SH_6 N_MM18_g 0.0010039f
cc_235 N_SH_14 N_CLKN_10 0.00226816f
cc_236 N_SH_5 N_MM12_g 0.00951832f
cc_237 N_SH_14 N_MM18_g 0.0162704f
cc_238 N_SH_5 N_CLKB_22 0.000127039f
cc_239 N_SH_6 N_MM13_g 0.000141727f
cc_240 N_SH_18 N_CLKB_19 0.000214844f
cc_241 N_SH_14 N_MM13_g 0.00675261f
cc_242 N_SH_13 N_MM13_g 0.00679213f
cc_243 N_SH_23 N_CLKB_19 0.000307038f
cc_244 N_SH_25 N_CLKB_19 0.000945889f
cc_245 N_SH_16 N_CLKB_2 0.000463902f
cc_246 N_SH_17 N_CLKB_19 0.000531726f
cc_247 N_SH_5 N_CLKB_2 0.000532303f
cc_248 N_SH_15 N_CLKB_19 0.000558577f
cc_249 N_SH_15 N_CLKB_22 0.00106396f
cc_250 N_SH_16 N_CLKB_19 0.00407655f
cc_251 N_SH_5 N_MM13_g 0.0184248f
cc_252 N_SH_16 N_NET029_3 0.00011607f
cc_253 N_SH_23 N_NET029_3 0.000158302f
cc_254 N_SH_14 N_NET029_3 0.000437544f
cc_255 N_SH_13 N_NET029_3 0.000465189f
cc_256 N_SH_6 N_NET029_4 0.000685919f
cc_257 N_SH_23 N_NET029_4 0.000294199f
cc_258 N_SH_23 N_NET029_17 0.000539863f
cc_259 N_SH_15 N_NET029_16 0.000589582f
cc_260 N_SH_14 N_NET029_4 0.000599882f
cc_261 N_SH_15 N_NET029_18 0.00168479f
cc_262 N_SH_5 N_NET029_3 0.00372999f
cc_263 N_SH_15 N_MM19_g 0.000112895f
cc_264 N_SH_17 N_MM19_g 0.000139439f
cc_265 N_SH_22 N_MM19_g 0.00019066f
cc_266 N_SH_27 N_MM19_g 0.000199208f
cc_267 N_SH_26 N_SS_12 0.000219151f
cc_268 N_MM14_g N_SS_10 0.00686366f
cc_269 N_MM14_g N_SS_11 0.00682864f
cc_270 N_SH_20 N_SS_4 0.000249533f
cc_271 N_SH_22 N_SS_15 0.00709845f
cc_272 N_SH_2 N_SS_15 0.00028578f
cc_273 N_SH_21 N_SS_15 0.00183608f
cc_274 N_MM14_g N_SS_3 0.000405f
cc_275 N_MM14_g N_SS_4 0.000527123f
cc_276 N_SH_20 N_SS_14 0.00065136f
cc_277 N_SH_1 N_SS_1 0.00070153f
cc_278 N_SH_24 N_SS_16 0.000793581f
cc_279 N_SH_16 N_SS_1 0.000844674f
cc_280 N_SH_27 N_SS_15 0.000900659f
cc_281 N_SH_19 N_SS_12 0.000953822f
cc_282 N_SH_21 N_SS_13 0.00105754f
cc_283 N_MM14_g N_SS_1 0.00110551f
cc_284 N_SH_1 N_MM19_g 0.00113663f
cc_285 N_SH_27 N_SS_14 0.00125874f
cc_286 N_SH_18 N_SS_12 0.00159032f
cc_287 N_SH_28 N_SS_15 0.00188796f
cc_288 N_SH_16 N_SS_12 0.00474118f
cc_289 N_MM14_g N_MM19_g 0.0294855f
x_PM_DFFLQNx1_ASAP7_75t_R%CLKN VSS N_MM22_g N_MM1_g N_MM9_g N_MM12_g N_MM18_g
+ N_MM20_d N_MM21_d N_CLKN_28 N_CLKN_35 N_CLKN_32 N_CLKN_9 N_CLKN_34 N_CLKN_8
+ N_CLKN_21 N_CLKN_22 N_CLKN_26 N_CLKN_25 N_CLKN_1 N_CLKN_27 N_CLKN_36
+ N_CLKN_23 N_CLKN_29 N_CLKN_2 N_CLKN_5 N_CLKN_30 N_CLKN_3 N_CLKN_10 N_CLKN_31
+ N_CLKN_33 N_CLKN_24 PM_DFFLQNx1_ASAP7_75t_R%CLKN
cc_290 N_CLKN_28 N_MM20_g 8.64818e-20
cc_291 N_CLKN_35 N_MM20_g 8.69563e-20
cc_292 N_CLKN_32 N_MM20_g 0.000192798f
cc_293 N_CLKN_9 N_MM20_g 0.00109915f
cc_294 N_CLKN_34 N_MM20_g 0.000233607f
cc_295 N_CLKN_8 N_MM20_g 0.00117509f
cc_296 N_CLKN_21 N_MM20_g 0.0112203f
cc_297 N_CLKN_22 N_MM20_g 0.0113257f
cc_298 N_CLKN_26 N_CLK_8 0.000734123f
cc_299 N_CLKN_25 N_CLK_5 0.000758513f
cc_300 N_CLKN_1 N_CLK_8 0.000777867f
cc_301 N_CLKN_27 N_CLK_1 0.000922771f
cc_302 N_CLKN_26 N_CLK_6 0.00131231f
cc_303 N_CLKN_27 N_CLK_7 0.00136564f
cc_304 N_CLKN_36 N_CLK_8 0.00169579f
cc_305 N_CLKN_23 N_CLK_4 0.00177586f
cc_306 N_CLKN_27 N_CLK_4 0.00214909f
cc_307 N_CLKN_34 N_CLK_8 0.00227131f
cc_308 N_CLKN_25 N_CLK_7 0.00227493f
cc_309 N_CLKN_1 N_CLK_1 0.00232584f
cc_310 N_CLKN_27 N_CLK_8 0.00241801f
cc_311 N_CLKN_32 N_CLK_8 0.00279116f
cc_312 N_MM22_g N_MM20_g 0.0351395f
*END of DFFLQNx1_ASAP7_75t_R.pxi
.ENDS
** Design:	DFFLQNx2_ASAP7_75t_R
* Created:	"Fri Aug 17 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "DFFLQNx2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "DFFLQNx2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_DFFLQNx2_ASAP7_75t_R%noxref_26 VSS 1
c1 1 VSS 0.0415127f
.ends

.subckt PM_DFFLQNx2_ASAP7_75t_R%noxref_29 VSS 1
c1 1 VSS 0.04235f
.ends

.subckt PM_DFFLQNx2_ASAP7_75t_R%noxref_28 VSS 1
c1 1 VSS 0.0423692f
.ends

.subckt PM_DFFLQNx2_ASAP7_75t_R%QN VSS 21 16 17 28 29 7 8 11 1 2
c1 1 VSS 0.0101807f
c2 2 VSS 0.0110509f
c3 7 VSS 0.00454138f
c4 8 VSS 0.00456959f
c5 9 VSS 0.00897496f
c6 10 VSS 0.00972674f
c7 11 VSS 0.00761679f
c8 12 VSS 0.00349085f
c9 13 VSS 0.00344944f
r1 29 27 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0430 $Y=0.2025 $X2=1.0405 $Y2=0.2025
r2 2 27 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0260 $Y=0.2025 $X2=1.0405 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0115 $Y=0.2025 $X2=1.0260 $Y2=0.2025
r4 28 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0090 $Y=0.2025 $X2=1.0115 $Y2=0.2025
r5 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0260 $Y=0.2025
+ $X2=1.0260 $Y2=0.2340
r6 24 25 9.32759 $w=1.3e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.2340 $X2=1.0660 $Y2=0.2340
r7 10 24 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.0145
+ $Y=0.2340 $X2=1.0260 $Y2=0.2340
r8 13 23 7.2121 $w=1.53211e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1060 $Y=0.2340 $X2=1.1060 $Y2=0.1960
r9 13 25 7.67848 $w=1.4125e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=1.1060
+ $Y=0.2340 $X2=1.0660 $Y2=0.2340
r10 22 23 9.73567 $w=1.3e-08 $l=4.18e-08 $layer=M1 $thickness=3.6e-08 $X=1.1060
+ $Y=0.1542 $X2=1.1060 $Y2=0.1960
r11 21 22 3.08976 $w=1.3e-08 $l=1.32e-08 $layer=M1 $thickness=3.6e-08 $X=1.1060
+ $Y=0.1410 $X2=1.1060 $Y2=0.1542
r12 21 20 6.00464 $w=1.3e-08 $l=2.58e-08 $layer=M1 $thickness=3.6e-08 $X=1.1060
+ $Y=0.1410 $X2=1.1060 $Y2=0.1152
r13 11 12 5.69636 $w=1.58e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1060 $Y=0.0675 $X2=1.1060 $Y2=0.0360
r14 11 20 11.1348 $w=1.3e-08 $l=4.77e-08 $layer=M1 $thickness=3.6e-08 $X=1.1060
+ $Y=0.0675 $X2=1.1060 $Y2=0.1152
r15 12 19 7.67848 $w=1.4125e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=1.1060
+ $Y=0.0360 $X2=1.0660 $Y2=0.0360
r16 18 19 9.32759 $w=1.3e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.0360 $X2=1.0660 $Y2=0.0360
r17 9 18 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.0145
+ $Y=0.0360 $X2=1.0260 $Y2=0.0360
r18 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0260 $Y=0.0675
+ $X2=1.0260 $Y2=0.0360
r19 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.0430 $Y=0.0675 $X2=1.0405 $Y2=0.0675
r20 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.0260 $Y=0.0675 $X2=1.0405 $Y2=0.0675
r21 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.0115 $Y=0.0675 $X2=1.0260 $Y2=0.0675
r22 16 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.0090 $Y=0.0675 $X2=1.0115 $Y2=0.0675
.ends

.subckt PM_DFFLQNx2_ASAP7_75t_R%noxref_27 VSS 1
c1 1 VSS 0.0415045f
.ends

.subckt PM_DFFLQNx2_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.00423603f
.ends

.subckt PM_DFFLQNx2_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.00433496f
.ends

.subckt PM_DFFLQNx2_ASAP7_75t_R%PD3 VSS 2 4 1
c1 1 VSS 0.000984951f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0405 $X2=0.4905 $Y2=0.0405
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0405 $X2=0.4735 $Y2=0.0405
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4735 $Y=0.0405 $X2=0.4905 $Y2=0.0405
.ends

.subckt PM_DFFLQNx2_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.00417384f
.ends

.subckt PM_DFFLQNx2_ASAP7_75t_R%PD4 VSS 2 4 1
c1 1 VSS 0.00094851f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.2295 $X2=0.7605 $Y2=0.2295
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.2295 $X2=0.7435 $Y2=0.2295
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7435 $Y=0.2295 $X2=0.7605 $Y2=0.2295
.ends

.subckt PM_DFFLQNx2_ASAP7_75t_R%PU1 VSS 2 4 1
c1 1 VSS 0.00097377f
r1 4 3 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3365 $Y2=0.2025
r2 2 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3195 $Y2=0.2025
r3 1 3 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3195 $Y=0.2025 $X2=0.3365 $Y2=0.2025
.ends

.subckt PM_DFFLQNx2_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.00418892f
.ends

.subckt PM_DFFLQNx2_ASAP7_75t_R%SS VSS 9 31 40 12 10 11 4 15 3 14 1 16 13
c1 1 VSS 0.00107529f
c2 3 VSS 0.00625572f
c3 4 VSS 0.00661474f
c4 9 VSS 0.0384302f
c5 10 VSS 0.00321469f
c6 11 VSS 0.00320919f
c7 12 VSS 0.00183356f
c8 13 VSS 0.0134807f
c9 14 VSS 0.00921502f
c10 15 VSS 0.00711838f
c11 16 VSS 0.00323752f
c12 17 VSS 0.0034663f
c13 18 VSS 0.00338942f
r1 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.2295 $X2=0.8620 $Y2=0.2295
r2 40 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.2295 $X2=0.8495 $Y2=0.2295
r3 4 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.2295
+ $X2=0.8640 $Y2=0.2340
r4 37 38 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.2340 $X2=0.8865 $Y2=0.2340
r5 14 18 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9180 $Y=0.2340 $X2=0.9450 $Y2=0.2340
r6 14 38 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.2340 $X2=0.8865 $Y2=0.2340
r7 18 35 6.74572 $w=1.545e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.2340 $X2=0.9450 $Y2=0.1980
r8 34 35 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1690 $X2=0.9450 $Y2=0.1980
r9 33 34 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1420 $X2=0.9450 $Y2=0.1690
r10 32 33 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1035 $X2=0.9450 $Y2=0.1420
r11 15 17 5.69636 $w=1.58e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.0675 $X2=0.9450 $Y2=0.0360
r12 15 32 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.0675 $X2=0.9450 $Y2=0.1035
r13 10 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.0405 $X2=0.8620 $Y2=0.0405
r14 31 10 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.0405 $X2=0.8495 $Y2=0.0405
r15 17 29 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.0360 $X2=0.9180 $Y2=0.0360
r16 3 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.0405
+ $X2=0.8640 $Y2=0.0360
r17 28 29 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.0360 $X2=0.9180 $Y2=0.0360
r18 27 28 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.0360 $X2=0.8910 $Y2=0.0360
r19 26 27 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.0360 $X2=0.8640 $Y2=0.0360
r20 13 16 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.0360 $X2=0.7830 $Y2=0.0360
r21 13 26 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0360 $X2=0.8370 $Y2=0.0360
r22 12 23 8.04505 $w=1.3e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.0705 $X2=0.7830 $Y2=0.1050
r23 12 16 6.39593 $w=1.55565e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7830 $Y=0.0705 $X2=0.7830 $Y2=0.0360
r24 1 20 2.36633 $w=2.3e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.7830
+ $Y=0.1055 $X2=0.7830 $Y2=0.1055
r25 1 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7830 $Y=0.1055
+ $X2=0.7830 $Y2=0.1050
r26 9 20 0.314665 $w=2.27e-07 $l=2.95e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.7830 $Y=0.1350 $X2=0.7830 $Y2=0.1055
.ends

.subckt PM_DFFLQNx2_ASAP7_75t_R%MS VSS 10 39 42 47 49 3 11 12 13 15 1 17 4 18
+ 14 16
c1 1 VSS 0.00219633f
c2 3 VSS 0.00537256f
c3 4 VSS 0.00935116f
c4 10 VSS 0.0374963f
c5 11 VSS 0.00285909f
c6 12 VSS 0.00269089f
c7 13 VSS 0.00225386f
c8 14 VSS 0.00186733f
c9 15 VSS 0.00403501f
c10 16 VSS 0.00298971f
c11 17 VSS 0.00101527f
c12 18 VSS 0.000434788f
c13 19 VSS 0.00295183f
r1 49 48 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.2295 $X2=0.6625 $Y2=0.2295
r2 13 48 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6500 $Y=0.2295 $X2=0.6625 $Y2=0.2295
r3 12 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2295 $X2=0.5920 $Y2=0.2295
r4 47 12 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.2295 $X2=0.5795 $Y2=0.2295
r5 44 13 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6210 $Y=0.2295 $X2=0.6480 $Y2=0.2295
r6 4 44 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08 $X=0.5940
+ $Y=0.2295 $X2=0.6210 $Y2=0.2295
r7 4 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2295
+ $X2=0.5965 $Y2=0.2340
r8 15 19 4.06404 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5965 $Y=0.2340 $X2=0.6210 $Y2=0.2340
r9 42 41 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.0405 $X2=0.6085 $Y2=0.0405
r10 40 41 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6040 $Y=0.0405 $X2=0.6085 $Y2=0.0405
r11 3 40 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5920 $Y=0.0405 $X2=0.6040 $Y2=0.0405
r12 11 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.0405 $X2=0.5920 $Y2=0.0405
r13 39 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0405 $X2=0.5795 $Y2=0.0405
r14 19 35 3.01468 $w=1.741e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.2340 $X2=0.6210 $Y2=0.2140
r15 3 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0405
+ $X2=0.5940 $Y2=0.0540
r16 34 35 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1850 $X2=0.6210 $Y2=0.2140
r17 33 34 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1660 $X2=0.6210 $Y2=0.1850
r18 32 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1525 $X2=0.6210 $Y2=0.1660
r19 31 32 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1310 $X2=0.6210 $Y2=0.1525
r20 17 28 3.60008 $w=1.51951e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.1105 $X2=0.6210 $Y2=0.0900
r21 17 31 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1105 $X2=0.6210 $Y2=0.1310
r22 16 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0540 $X2=0.5940 $Y2=0.0720
r23 27 28 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6075 $Y=0.0900 $X2=0.6210 $Y2=0.0900
r24 18 26 1.38478 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5940 $Y=0.0900 $X2=0.5830 $Y2=0.0900
r25 18 27 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5940 $Y=0.0900 $X2=0.6075 $Y2=0.0900
r26 18 29 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0900 $X2=0.5940 $Y2=0.0720
r27 25 26 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5515
+ $Y=0.0900 $X2=0.5830 $Y2=0.0900
r28 24 25 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0900 $X2=0.5515 $Y2=0.0900
r29 14 24 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5000
+ $Y=0.0900 $X2=0.5130 $Y2=0.0900
r30 1 21 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.5130
+ $Y=0.0900 $X2=0.5130 $Y2=0.0900
r31 1 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.0900
+ $X2=0.5130 $Y2=0.0900
r32 10 21 0.314665 $w=2.27e-07 $l=4.5e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5130 $Y2=0.0900
.ends

.subckt PM_DFFLQNx2_ASAP7_75t_R%PD2 VSS 7 12 5 1 4
c1 1 VSS 0.00727636f
c2 4 VSS 0.00188706f
c3 5 VSS 0.00233436f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4880 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r3 9 5 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.4605
+ $Y=0.2295 $X2=0.4860 $Y2=0.2295
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.4455
+ $Y=0.2295 $X2=0.4605 $Y2=0.2295
r5 1 8 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4320
+ $Y=0.2295 $X2=0.4455 $Y2=0.2295
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2295 $X2=0.4300 $Y2=0.2295
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2295 $X2=0.4175 $Y2=0.2295
.ends

.subckt PM_DFFLQNx2_ASAP7_75t_R%PD5 VSS 7 12 1 4 5
c1 1 VSS 0.0074664f
c2 4 VSS 0.00187629f
c3 5 VSS 0.00237792f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.0405 $X2=0.7705 $Y2=0.0405
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7580 $Y=0.0405 $X2=0.7705 $Y2=0.0405
r3 9 5 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.7425
+ $Y=0.0405 $X2=0.7560 $Y2=0.0405
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.7275
+ $Y=0.0405 $X2=0.7425 $Y2=0.0405
r5 1 8 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.7020
+ $Y=0.0405 $X2=0.7275 $Y2=0.0405
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.0405 $X2=0.7000 $Y2=0.0405
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.0405 $X2=0.6875 $Y2=0.0405
.ends

.subckt PM_DFFLQNx2_ASAP7_75t_R%PD1 VSS 7 10 5 4 1
c1 1 VSS 0.00972744f
c2 4 VSS 0.00316965f
c3 5 VSS 0.00186048f
r1 10 9 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r2 8 9 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r3 5 8 0.123457 $w=8.1e-08 $l=1e-08 $layer=N_src_drn $thickness=1e-09 $X=0.3780
+ $Y=0.0675 $X2=0.3880 $Y2=0.0675
r4 4 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3220 $Y2=0.0675
r5 7 4 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r6 1 5 1e-05
.ends

.subckt PM_DFFLQNx2_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.00478752f
.ends

.subckt PM_DFFLQNx2_ASAP7_75t_R%D VSS 9 3 4 1 6 5
c1 1 VSS 0.00681582f
c2 3 VSS 0.0834271f
c3 4 VSS 0.00585828f
c4 5 VSS 0.0068338f
c5 6 VSS 0.00763261f
r1 6 13 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.2340 $X2=0.2970 $Y2=0.2140
r2 5 8 5.17411 $w=1.46514e-08 $l=2.72e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0360 $X2=0.2970 $Y2=0.0632
r3 12 13 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1735 $X2=0.2970 $Y2=0.2140
r4 11 12 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1735
r5 9 10 2.85657 $w=1.3e-08 $l=1.22e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0820 $X2=0.2970 $Y2=0.0942
r6 9 8 4.37231 $w=1.3e-08 $l=1.88e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0820 $X2=0.2970 $Y2=0.0632
r7 4 10 5.07188 $w=1.3e-08 $l=2.18e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1160 $X2=0.2970 $Y2=0.0942
r8 4 11 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1160 $X2=0.2970 $Y2=0.1350
r9 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r10 1 11 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_DFFLQNx2_ASAP7_75t_R%SH VSS 11 12 13 70 73 77 80 16 24 26 14 6 19 17
+ 18 15 5 29 2 23 28 27 21 22 1 25 20
c1 1 VSS 0.000665047f
c2 2 VSS 0.00845479f
c3 5 VSS 0.00476783f
c4 6 VSS 0.00537673f
c5 11 VSS 0.0374716f
c6 12 VSS 0.0809929f
c7 13 VSS 0.080766f
c8 14 VSS 0.00519645f
c9 15 VSS 0.00537376f
c10 16 VSS 0.00849956f
c11 17 VSS 0.00207809f
c12 18 VSS 0.0018946f
c13 19 VSS 0.00280361f
c14 20 VSS 0.000861472f
c15 21 VSS 0.000540199f
c16 22 VSS 0.00135425f
c17 23 VSS 0.00399346f
c18 24 VSS 0.00614582f
c19 25 VSS 0.00231538f
c20 26 VSS 0.000137504f
c21 27 VSS 0.000413455f
c22 28 VSS 0.000388944f
c23 29 VSS 0.0116813f
r1 80 79 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r2 5 79 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6500 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r3 76 5 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6380 $Y=0.0405 $X2=0.6500 $Y2=0.0405
r4 14 76 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0405 $X2=0.6380 $Y2=0.0405
r5 77 14 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.0405 $X2=0.6335 $Y2=0.0405
r6 13 65 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=1.0530
+ $Y=0.1350 $X2=1.0530 $Y2=0.1350
r7 12 57 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.9990 $Y=0.1350 $X2=0.9990 $Y2=0.1350
r8 73 72 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r9 71 72 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7120 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r10 6 71 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7000 $Y=0.2295 $X2=0.7120 $Y2=0.2295
r11 15 6 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.2295 $X2=0.7000 $Y2=0.2295
r12 70 15 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.2295 $X2=0.6875 $Y2=0.2295
r13 5 55 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.0405
+ $X2=0.6480 $Y2=0.0360
r14 63 65 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.0405 $Y=0.1350 $X2=1.0530 $Y2=0.1350
r15 62 63 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.0260 $Y=0.1350 $X2=1.0405 $Y2=0.1350
r16 60 62 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.0115 $Y=0.1350 $X2=1.0260 $Y2=0.1350
r17 58 60 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=1.0085 $Y=0.1350 $X2=1.0115 $Y2=0.1350
r18 57 58 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.9990
+ $Y=0.1350 $X2=1.0085 $Y2=0.1350
r19 2 57 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.9895
+ $Y=0.1350 $X2=0.9990 $Y2=0.1350
r20 6 48 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7020 $Y=0.2295
+ $X2=0.7020 $Y2=0.2340
r21 55 56 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6480
+ $Y=0.0360 $X2=0.6615 $Y2=0.0360
r22 53 56 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0360 $X2=0.6615 $Y2=0.0360
r23 52 53 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6860
+ $Y=0.0360 $X2=0.6750 $Y2=0.0360
r24 16 25 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.7040
+ $Y=0.0360 $X2=0.7290 $Y2=0.0360
r25 16 52 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7040
+ $Y=0.0360 $X2=0.6860 $Y2=0.0360
r26 50 57 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.9990 $Y=0.1440
+ $X2=0.9990 $Y2=0.1350
r27 23 50 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.9990
+ $Y=0.1080 $X2=0.9990 $Y2=0.1440
r28 48 49 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.2340 $X2=0.7155 $Y2=0.2340
r29 24 49 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.2340 $X2=0.7155 $Y2=0.2340
r30 25 41 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.0360 $X2=0.7290 $Y2=0.0630
r31 45 50 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.9990 $Y=0.1530
+ $X2=0.9990 $Y2=0.1440
r32 44 45 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1530 $X2=0.9990 $Y2=0.1530
r33 43 44 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1530 $X2=0.9450 $Y2=0.1530
r34 29 43 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.8795
+ $Y=0.1530 $X2=0.8910 $Y2=0.1530
r35 42 43 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.8910 $Y=0.1485 $X2=0.8910
+ $Y2=0.1530
r36 22 42 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1305 $X2=0.8910 $Y2=0.1485
r37 18 37 6.50021 $w=1.33448e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1980 $X2=0.7290 $Y2=0.1690
r38 18 24 7.21452 $w=1.425e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1980 $X2=0.7290 $Y2=0.2340
r39 40 41 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.0900 $X2=0.7290 $Y2=0.0630
r40 39 40 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1090 $X2=0.7290 $Y2=0.0900
r41 17 26 4.67854 $w=1.44583e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1360 $X2=0.7290 $Y2=0.1600
r42 17 39 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1360 $X2=0.7290 $Y2=0.1090
r43 28 38 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1575 $X2=0.8910 $Y2=0.1665
r44 28 42 1.50855 $w=1.55e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1575 $X2=0.8910 $Y2=0.1485
r45 28 43 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.8910 $Y=0.1575 $X2=0.8910
+ $Y2=0.1530
r46 26 37 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1600 $X2=0.7290 $Y2=0.1690
r47 36 38 4.19024 $w=1.156e-08 $l=2.54018e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8660 $Y=0.1620 $X2=0.8910 $Y2=0.1665
r48 21 27 1.38478 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8480 $Y=0.1620 $X2=0.8370 $Y2=0.1620
r49 21 36 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8480
+ $Y=0.1620 $X2=0.8660 $Y2=0.1620
r50 35 37 4.4015 $w=1.35e-08 $l=2.78927e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7560 $Y=0.1620 $X2=0.7290 $Y2=0.1690
r51 34 35 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1620 $X2=0.7560 $Y2=0.1620
r52 19 27 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.1620 $X2=0.8370 $Y2=0.1620
r53 19 34 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.1620 $X2=0.7830 $Y2=0.1620
r54 27 33 4.88263 $w=1.47308e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8370 $Y=0.1620 $X2=0.8370 $Y2=0.1360
r55 20 33 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1180 $X2=0.8370 $Y2=0.1360
r56 11 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.8370
+ $Y=0.1350 $X2=0.8370 $Y2=0.1350
r57 1 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8370 $Y=0.1350
+ $X2=0.8370 $Y2=0.1360
.ends

.subckt PM_DFFLQNx2_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.00469434f
.ends

.subckt PM_DFFLQNx2_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.0418056f
.ends

.subckt PM_DFFLQNx2_ASAP7_75t_R%CLK VSS 11 3 8 5 1 6 7 4
c1 1 VSS 0.00262062f
c2 3 VSS 0.0598043f
c3 4 VSS 0.00105427f
c4 5 VSS 0.00414517f
c5 6 VSS 0.00373949f
c6 7 VSS 0.00235261f
c7 8 VSS 0.00199015f
r1 6 17 3.22357 $w=2.26279e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.2125 $X2=0.1080 $Y2=0.1820
r2 5 15 3.22357 $w=2.26279e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0575 $X2=0.1080 $Y2=0.0880
r3 16 17 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.1820 $X2=0.1080 $Y2=0.1820
r4 8 13 2.6406 $w=2.38947e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1820 $X2=0.0810 $Y2=0.1540
r5 8 16 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1820 $X2=0.0945 $Y2=0.1820
r6 14 15 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.0880 $X2=0.1080 $Y2=0.0880
r7 7 10 1.76614 $w=2.65738e-08 $l=2.42e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0880 $X2=0.0810 $Y2=0.1122
r8 7 14 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0880 $X2=0.0945 $Y2=0.0880
r9 11 12 0.874462 $w=1.3e-08 $l=3.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1227
r10 11 10 1.57403 $w=1.3e-08 $l=6.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1122
r11 4 12 2.85657 $w=1.3e-08 $l=1.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1227
r12 4 13 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1540
r13 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r14 1 4 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_DFFLQNx2_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.0418511f
.ends

.subckt PM_DFFLQNx2_ASAP7_75t_R%MH VSS 9 47 51 57 61 10 20 3 16 1 17 4 12 14 18
+ 15 19
c1 1 VSS 0.0002757f
c2 3 VSS 0.00624436f
c3 4 VSS 0.00540897f
c4 9 VSS 0.0364051f
c5 10 VSS 0.0022711f
c6 11 VSS 9.01122e-20
c7 12 VSS 0.00278109f
c8 13 VSS 6.89826e-20
c9 14 VSS 0.00852254f
c10 15 VSS 0.00125695f
c11 16 VSS 0.000667797f
c12 17 VSS 0.000550194f
c13 18 VSS 0.00649713f
c14 19 VSS 1.21302e-20
c15 20 VSS 0.00228322f
r1 61 60 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r2 59 60 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r3 3 59 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3760 $Y=0.2295 $X2=0.3880 $Y2=0.2295
r4 13 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2295 $X2=0.3760 $Y2=0.2295
r5 55 56 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r6 57 55 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.1890 $X2=0.3635 $Y2=0.1890
r7 12 56 0.185185 $w=5.4e-08 $l=1e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r8 12 3 0.518519 $w=3.9e-08 $l=4.05494e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.1890 $X2=0.3760 $Y2=0.2295
r9 3 44 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2295
+ $X2=0.3780 $Y2=0.2340
r10 51 50 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r11 49 50 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4420 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r12 4 49 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4300 $Y=0.0405 $X2=0.4420 $Y2=0.0405
r13 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0405 $X2=0.4300 $Y2=0.0405
r14 10 4 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0810 $X2=0.4300 $Y2=0.0810
r15 47 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0810 $X2=0.4175 $Y2=0.0810
r16 44 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r17 42 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r18 41 42 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4160
+ $Y=0.2340 $X2=0.4050 $Y2=0.2340
r19 14 20 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4340
+ $Y=0.2340 $X2=0.4590 $Y2=0.2340
r20 14 41 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4340
+ $Y=0.2340 $X2=0.4160 $Y2=0.2340
r21 4 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0405
+ $X2=0.4320 $Y2=0.0360
r22 20 34 3.01468 $w=1.741e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4590 $Y2=0.2140
r23 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4455 $Y2=0.0360
r24 18 31 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4590 $Y2=0.0630
r25 18 37 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4455 $Y2=0.0360
r26 33 34 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1850 $X2=0.4590 $Y2=0.2140
r27 32 33 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1660 $X2=0.4590 $Y2=0.1850
r28 16 19 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1525 $X2=0.4590 $Y2=0.1310
r29 16 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1525 $X2=0.4590 $Y2=0.1660
r30 30 31 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0900 $X2=0.4590 $Y2=0.0630
r31 29 30 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1025 $X2=0.4590 $Y2=0.0900
r32 15 19 2.78392 $w=1.56471e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1140 $X2=0.4590 $Y2=0.1310
r33 15 29 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1140 $X2=0.4590 $Y2=0.1025
r34 19 27 4.18306 $w=1.49565e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1310 $X2=0.4820 $Y2=0.1310
r35 26 27 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5000
+ $Y=0.1310 $X2=0.4820 $Y2=0.1310
r36 25 26 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1310 $X2=0.5000 $Y2=0.1310
r37 17 24 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1310 $X2=0.5670 $Y2=0.1310
r38 17 25 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1310 $X2=0.5130 $Y2=0.1310
r39 23 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1330
+ $X2=0.5670 $Y2=0.1310
r40 1 22 1.47681 $w=1.53e-08 $l=9e-09 $layer=LIG $thickness=4.8e-08 $X=0.5670
+ $Y=0.1215 $X2=0.5670 $Y2=0.1305
r41 22 23 5.31651 $w=1.53e-08 $l=2.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.5670 $Y=0.1305 $X2=0.5670 $Y2=0.1330
r42 9 22 0.314665 $w=2.27e-07 $l=4.5e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5670 $Y=0.1350 $X2=0.5670 $Y2=0.1305
r43 3 12 1e-05
.ends

.subckt PM_DFFLQNx2_ASAP7_75t_R%CLKN VSS 16 17 18 19 20 99 101 28 35 32 9 34 8
+ 21 22 26 25 1 27 36 23 29 2 5 30 3 10 31 33 24
c1 1 VSS 0.00148346f
c2 2 VSS 0.000298605f
c3 3 VSS 7.25213e-20
c4 4 VSS 1e-36
c5 5 VSS 0.000425464f
c6 8 VSS 0.00771357f
c7 9 VSS 0.00771771f
c8 10 VSS 0.0035511f
c9 16 VSS 0.0590851f
c10 17 VSS 0.00561042f
c11 18 VSS 0.00511489f
c12 19 VSS 0.00438046f
c13 20 VSS 0.00517375f
c14 21 VSS 0.00655992f
c15 22 VSS 0.00651045f
c16 23 VSS 0.00804227f
c17 24 VSS 0.00180784f
c18 25 VSS 0.00454209f
c19 26 VSS 0.00375644f
c20 27 VSS 0.000658467f
c21 28 VSS 0.000261285f
c22 29 VSS 0.000827042f
c23 30 VSS 0.00146342f
c24 31 VSS 0.00383266f
c25 32 VSS 0.00190647f
c26 33 VSS 0.00393343f
c27 34 VSS 0.00084146f
c28 35 VSS 0.000477398f
c29 36 VSS 0.0228768f
r1 101 100 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r2 22 100 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r3 99 98 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r4 21 98 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r5 9 96 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0550 $Y2=0.2340
r6 8 93 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0550 $Y2=0.0360
r7 95 96 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.2340 $X2=0.0550 $Y2=0.2340
r8 26 95 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0460 $Y2=0.2340
r9 26 33 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0180 $Y2=0.2340
r10 92 93 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.0360 $X2=0.0550 $Y2=0.0360
r11 25 92 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0460 $Y2=0.0360
r12 25 31 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0180 $Y2=0.0360
r13 5 91 2.78395 $w=2.4e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08 $X=0.7290
+ $Y=0.1780 $X2=0.7250 $Y2=0.1780
r14 20 5 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.7290 $Y=0.1350 $X2=0.7290 $Y2=0.1780
r15 4 84 10.3807 $w=2.30357e-08 $l=0 $layer=LISD $thickness=3.675e-08 $X=0.6210
+ $Y=0.1780 $X2=0.6210 $Y2=0.1780
r16 19 4 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.6210 $Y=0.1350 $X2=0.6210 $Y2=0.1780
r17 3 77 2.78395 $w=2.4e-08 $l=5e-09 $layer=LIG $thickness=4.8e-08 $X=0.4590
+ $Y=0.1780 $X2=0.4640 $Y2=0.1780
r18 18 3 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4590 $Y2=0.1780
r19 33 72 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.2340 $X2=0.0180 $Y2=0.2125
r20 31 71 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.0360 $X2=0.0180 $Y2=0.0575
r21 90 91 4.8113 $w=2.22e-08 $l=1.5e-09 $layer=LISD $thickness=2.7e-08
+ $X=0.7235 $Y=0.1780 $X2=0.7250 $Y2=0.1780
r22 89 90 10.8887 $w=2.22e-08 $l=2.15e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7020 $Y=0.1780 $X2=0.7235 $Y2=0.1780
r23 88 89 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6885 $Y=0.1780 $X2=0.7020 $Y2=0.1780
r24 87 88 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6750 $Y=0.1780 $X2=0.6885 $Y2=0.1780
r25 86 87 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6615 $Y=0.1780 $X2=0.6750 $Y2=0.1780
r26 85 86 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6480 $Y=0.1780 $X2=0.6615 $Y2=0.1780
r27 84 85 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6210 $Y=0.1780 $X2=0.6480 $Y2=0.1780
r28 83 84 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5940 $Y=0.1780 $X2=0.6210 $Y2=0.1780
r29 82 83 7.09034 $w=2.22e-08 $l=1.4e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5800 $Y=0.1780 $X2=0.5940 $Y2=0.1780
r30 81 82 6.58388 $w=2.22e-08 $l=1.3e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5670 $Y=0.1780 $X2=0.5800 $Y2=0.1780
r31 80 81 6.58388 $w=2.22e-08 $l=1.3e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5540 $Y=0.1780 $X2=0.5670 $Y2=0.1780
r32 79 80 7.09034 $w=2.22e-08 $l=1.4e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5400 $Y=0.1780 $X2=0.5540 $Y2=0.1780
r33 78 79 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5265 $Y=0.1780 $X2=0.5400 $Y2=0.1780
r34 76 77 10.3823 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4775 $Y=0.1780 $X2=0.4640 $Y2=0.1780
r35 75 76 11.142 $w=2.22e-08 $l=2.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4995 $Y=0.1780 $X2=0.4775 $Y2=0.1780
r36 74 78 1.51936 $w=2.22e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.5235
+ $Y=0.1780 $X2=0.5265 $Y2=0.1780
r37 73 74 5.31775 $w=2.22e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5130 $Y=0.1780 $X2=0.5235 $Y2=0.1780
r38 10 73 5.31775 $w=2.22e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5025 $Y=0.1780 $X2=0.5130 $Y2=0.1780
r39 10 75 1.51936 $w=2.22e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.5025
+ $Y=0.1780 $X2=0.4995 $Y2=0.1780
r40 2 65 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
r41 17 2 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r42 24 32 0.998523 $w=1.74118e-08 $l=1.01119e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1990 $X2=0.0165 $Y2=0.1890
r43 24 72 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1990 $X2=0.0180 $Y2=0.2125
r44 70 71 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0880 $X2=0.0180 $Y2=0.0575
r45 69 70 10.9599 $w=1.3e-08 $l=4.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1350 $X2=0.0180 $Y2=0.0880
r46 23 32 2.63085 $w=1.54194e-08 $l=1.7066e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1720 $X2=0.0165 $Y2=0.1890
r47 23 69 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1720 $X2=0.0180 $Y2=0.1350
r48 67 73 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5130 $Y=0.1845
+ $X2=0.5130 $Y2=0.1780
r49 30 67 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1680 $X2=0.5130 $Y2=0.1845
r50 65 66 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1555
r51 29 63 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1735 $X2=0.3510 $Y2=0.1890
r52 29 66 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1735 $X2=0.3510 $Y2=0.1555
r53 60 61 1.90199 $w=1.38333e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.0255 $Y=0.1890 $X2=0.0345 $Y2=0.1890
r54 32 60 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0165
+ $Y=0.1890 $X2=0.0255 $Y2=0.1890
r55 58 67 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.5130 $Y=0.1890
+ $X2=0.5130 $Y2=0.1845
r56 57 58 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.4320
+ $Y=0.1890 $X2=0.5130 $Y2=0.1890
r57 56 57 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1890 $X2=0.4320 $Y2=0.1890
r58 56 63 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.3510 $Y=0.1890
+ $X2=0.3510 $Y2=0.1890
r59 55 56 15.2739 $w=1.3e-08 $l=6.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.2855
+ $Y=0.1890 $X2=0.3510 $Y2=0.1890
r60 54 55 20.2875 $w=1.3e-08 $l=8.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.1985
+ $Y=0.1890 $X2=0.2855 $Y2=0.1890
r61 53 54 9.211 $w=1.3e-08 $l=3.95e-08 $layer=M2 $thickness=3.6e-08 $X=0.1590
+ $Y=0.1890 $X2=0.1985 $Y2=0.1890
r62 52 53 14.691 $w=1.3e-08 $l=6.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.0960
+ $Y=0.1890 $X2=0.1590 $Y2=0.1890
r63 51 52 14.691 $w=1.3e-08 $l=6.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.0330
+ $Y=0.1890 $X2=0.0960 $Y2=0.1890
r64 51 61 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.0330 $Y=0.1890
+ $X2=0.0345 $Y2=0.1890
r65 36 51 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.0215
+ $Y=0.1890 $X2=0.0330 $Y2=0.1890
r66 48 49 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1590
+ $Y=0.1890 $X2=0.1740 $Y2=0.1890
r67 48 53 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1590 $Y=0.1890
+ $X2=0.1590 $Y2=0.1890
r68 34 46 2.78392 $w=1.56471e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1890 $X2=0.1890 $Y2=0.1720
r69 34 49 2.31754 $w=1.6e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1890 $X2=0.1740 $Y2=0.1890
r70 28 35 2.78149 $w=1.76421e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1540 $X2=0.1890 $Y2=0.1350
r71 28 46 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1540 $X2=0.1890 $Y2=0.1720
r72 35 45 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1640 $Y2=0.1350
r73 44 45 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.1465
+ $Y=0.1350 $X2=0.1640 $Y2=0.1350
r74 43 44 0.46638 $w=1.3e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.1445
+ $Y=0.1350 $X2=0.1465 $Y2=0.1350
r75 42 43 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1445 $Y2=0.1350
r76 27 42 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1235
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r77 16 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r78 1 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
r79 9 22 1e-05
r80 8 21 1e-05
.ends

.subckt PM_DFFLQNx2_ASAP7_75t_R%CLKB VSS 11 12 57 59 17 6 5 16 15 13 21 22 14
+ 19 18 2 1 20
c1 1 VSS 4.22509e-20
c2 2 VSS 0.000150034f
c3 5 VSS 0.00727931f
c4 6 VSS 0.00729125f
c5 11 VSS 0.00437566f
c6 12 VSS 0.0045835f
c7 13 VSS 0.00646428f
c8 14 VSS 0.00647226f
c9 15 VSS 0.00858574f
c10 16 VSS 0.00855551f
c11 17 VSS 0.00621647f
c12 18 VSS 0.000545167f
c13 19 VSS 0.0015389f
c14 20 VSS 0.00360961f
c15 21 VSS 0.00300542f
c16 22 VSS 0.0162898f
r1 14 6 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1600 $Y2=0.2160
r2 59 14 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r3 13 5 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1600 $Y2=0.0540
r4 57 13 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r5 6 53 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r6 5 50 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r7 53 54 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1845 $Y2=0.2340
r8 16 21 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.2340 $X2=0.2430 $Y2=0.2340
r9 16 54 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.1845 $Y2=0.2340
r10 50 51 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1845 $Y2=0.0360
r11 15 20 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.0360 $X2=0.2430 $Y2=0.0360
r12 15 51 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.1845 $Y2=0.0360
r13 2 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6750 $Y=0.1350
+ $X2=0.6750 $Y2=0.1440
r14 12 2 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6750
+ $Y=0.1350 $X2=0.6750 $Y2=0.1350
r15 21 44 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.2340 $X2=0.2430 $Y2=0.2125
r16 20 41 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0360 $X2=0.2430 $Y2=0.0575
r17 19 45 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1125 $X2=0.6750 $Y2=0.1440
r18 43 44 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1990 $X2=0.2430 $Y2=0.2125
r19 42 43 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1890 $X2=0.2430 $Y2=0.1990
r20 40 41 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0880 $X2=0.2430 $Y2=0.0575
r21 39 40 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1160 $X2=0.2430 $Y2=0.0880
r22 38 42 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1710 $X2=0.2430 $Y2=0.1890
r23 37 38 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1530 $X2=0.2430 $Y2=0.1710
r24 17 37 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1530
r25 17 39 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1160
r26 35 45 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.6750 $Y=0.1530
+ $X2=0.6750 $Y2=0.1440
r27 34 35 18.3054 $w=1.3e-08 $l=7.85e-08 $layer=M2 $thickness=3.6e-08 $X=0.5965
+ $Y=0.1530 $X2=0.6750 $Y2=0.1530
r28 33 34 29.3819 $w=1.3e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.4705
+ $Y=0.1530 $X2=0.5965 $Y2=0.1530
r29 32 33 15.2739 $w=1.3e-08 $l=6.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1530 $X2=0.4705 $Y2=0.1530
r30 31 32 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1530 $X2=0.4050 $Y2=0.1530
r31 30 31 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1530 $X2=0.3240 $Y2=0.1530
r32 30 37 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.2430 $Y=0.1530
+ $X2=0.2430 $Y2=0.1530
r33 22 30 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.2315
+ $Y=0.1530 $X2=0.2430 $Y2=0.1530
r34 28 32 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4050 $Y=0.1440
+ $X2=0.4050 $Y2=0.1530
r35 18 28 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1160 $X2=0.4050 $Y2=0.1440
r36 11 1 5.63117 $w=1.26721e-07 $l=2e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4050 $Y2=0.1330
r37 1 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1330
+ $X2=0.4050 $Y2=0.1440
.ends


*
.SUBCKT DFFLQNx2_ASAP7_75t_R VSS VDD CLK D QN
*
* VSS VSS
* VDD VDD
* CLK CLK
* D D
* QN QN
*
*

MM20 N_MM20_d N_MM20_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM23 N_MM23_d N_MM22_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM10_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM6 N_MM6_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM12 N_MM12_d N_MM12_g N_MM12_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM17 N_MM17_d N_MM13_g N_MM17_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM16 N_MM16_d N_MM19_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM14 N_MM14_d N_MM14_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM24 N_MM24_d N_MM24_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@2 N_MM24@2_d N_MM24@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM21 N_MM21_d N_MM20_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM22 N_MM22_d N_MM22_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM13 N_MM13_d N_MM13_g N_MM13_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM18 N_MM18_d N_MM18_g N_MM18_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM19 N_MM19_d N_MM19_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM15 N_MM15_d N_MM14_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM25 N_MM25_d N_MM24_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@2 N_MM25@2_d N_MM24@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "DFFLQNx2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "DFFLQNx2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_DFFLQNx2_ASAP7_75t_R%noxref_26 VSS N_noxref_26_1
+ PM_DFFLQNx2_ASAP7_75t_R%noxref_26
cc_1 N_noxref_26_1 N_SS_10 0.000639876f
cc_2 N_noxref_26_1 N_MM24_g 0.00170854f
cc_3 N_noxref_26_1 N_noxref_24_1 0.00777053f
cc_4 N_noxref_26_1 N_noxref_25_1 0.000476655f
x_PM_DFFLQNx2_ASAP7_75t_R%noxref_29 VSS N_noxref_29_1
+ PM_DFFLQNx2_ASAP7_75t_R%noxref_29
cc_5 N_noxref_29_1 N_MM24@2_g 0.00146705f
cc_6 N_noxref_29_1 N_QN_8 0.000820572f
cc_7 N_noxref_29_1 N_noxref_28_1 0.00176908f
x_PM_DFFLQNx2_ASAP7_75t_R%noxref_28 VSS N_noxref_28_1
+ PM_DFFLQNx2_ASAP7_75t_R%noxref_28
cc_8 N_noxref_28_1 N_MM24@2_g 0.00146411f
cc_9 N_noxref_28_1 N_QN_7 0.000829388f
x_PM_DFFLQNx2_ASAP7_75t_R%QN VSS QN N_MM24_d N_MM24@2_d N_MM25_d N_MM25@2_d
+ N_QN_7 N_QN_8 N_QN_11 N_QN_1 N_QN_2 PM_DFFLQNx2_ASAP7_75t_R%QN
cc_10 N_QN_7 N_SH_23 0.00133782f
cc_11 N_QN_7 N_SH_2 0.000492032f
cc_12 N_QN_7 N_SH_29 0.00072955f
cc_13 N_QN_8 N_MM24@2_g 0.0307893f
cc_14 N_QN_11 N_SH_2 0.0012524f
cc_15 N_QN_1 N_SH_23 0.0016689f
cc_16 N_QN_2 N_MM24@2_g 0.00211994f
cc_17 N_QN_1 N_MM24@2_g 0.00217625f
cc_18 N_QN_8 N_SH_2 0.00476758f
cc_19 N_QN_7 N_MM24_g 0.0371716f
cc_20 N_QN_7 N_MM24@2_g 0.0682669f
x_PM_DFFLQNx2_ASAP7_75t_R%noxref_27 VSS N_noxref_27_1
+ PM_DFFLQNx2_ASAP7_75t_R%noxref_27
cc_21 N_noxref_27_1 N_SS_11 0.000627018f
cc_22 N_noxref_27_1 N_MM24_g 0.00172435f
cc_23 N_noxref_27_1 N_noxref_24_1 0.000478522f
cc_24 N_noxref_27_1 N_noxref_25_1 0.00776006f
cc_25 N_noxref_27_1 N_noxref_26_1 0.00124076f
x_PM_DFFLQNx2_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_DFFLQNx2_ASAP7_75t_R%noxref_24
cc_26 N_noxref_24_1 N_SS_10 0.0170381f
cc_27 N_noxref_24_1 N_SH_1 0.00018406f
cc_28 N_noxref_24_1 N_MM14_g 0.00593747f
x_PM_DFFLQNx2_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_DFFLQNx2_ASAP7_75t_R%noxref_25
cc_29 N_noxref_25_1 N_SS_11 0.0168784f
cc_30 N_noxref_25_1 N_SH_1 0.000168104f
cc_31 N_noxref_25_1 N_MM14_g 0.00602616f
cc_32 N_noxref_25_1 N_noxref_24_1 0.00153921f
x_PM_DFFLQNx2_ASAP7_75t_R%PD3 VSS N_MM9_s N_MM8_d N_PD3_1
+ PM_DFFLQNx2_ASAP7_75t_R%PD3
cc_33 N_PD3_1 N_MM9_g 0.00772306f
cc_34 N_PD3_1 N_MM11_g 0.00772858f
x_PM_DFFLQNx2_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_DFFLQNx2_ASAP7_75t_R%noxref_19
cc_35 N_noxref_19_1 N_MM20_g 0.00367453f
cc_36 N_noxref_19_1 N_CLKN_8 4.38676e-20
cc_37 N_noxref_19_1 N_CLKN_33 5.38656e-20
cc_38 N_noxref_19_1 N_CLKN_24 8.26328e-20
cc_39 N_noxref_19_1 N_CLKN_32 8.8491e-20
cc_40 N_noxref_19_1 N_CLKN_23 0.00027147f
cc_41 N_noxref_19_1 N_CLKN_9 0.00050327f
cc_42 N_noxref_19_1 N_CLKN_22 0.0277397f
cc_43 N_noxref_19_1 N_noxref_18_1 0.00204488f
x_PM_DFFLQNx2_ASAP7_75t_R%PD4 VSS N_MM18_s N_MM19_d N_PD4_1
+ PM_DFFLQNx2_ASAP7_75t_R%PD4
cc_44 N_PD4_1 N_MM18_g 0.00773055f
cc_45 N_PD4_1 N_MM19_g 0.00776247f
x_PM_DFFLQNx2_ASAP7_75t_R%PU1 VSS N_MM3_d N_MM1_s N_PU1_1
+ PM_DFFLQNx2_ASAP7_75t_R%PU1
cc_46 N_PU1_1 N_MM1_g 0.0169384f
cc_47 N_PU1_1 N_MM3_g 0.0170114f
x_PM_DFFLQNx2_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_DFFLQNx2_ASAP7_75t_R%noxref_18
cc_48 N_noxref_18_1 N_MM20_g 0.00369069f
cc_49 N_noxref_18_1 N_CLKN_8 0.000543714f
cc_50 N_noxref_18_1 N_CLKN_9 4.21487e-20
cc_51 N_noxref_18_1 N_CLKN_31 5.87318e-20
cc_52 N_noxref_18_1 N_CLKN_23 0.00038388f
cc_53 N_noxref_18_1 N_CLKN_21 0.0276347f
x_PM_DFFLQNx2_ASAP7_75t_R%SS VSS N_MM19_g N_MM14_d N_MM15_d N_SS_12 N_SS_10
+ N_SS_11 N_SS_4 N_SS_15 N_SS_3 N_SS_14 N_SS_1 N_SS_16 N_SS_13
+ PM_DFFLQNx2_ASAP7_75t_R%SS
cc_54 N_MM19_g N_CLKN_10 0.000218803f
cc_55 N_MM19_g N_CLKN_5 0.000537557f
cc_56 N_MM19_g N_MM18_g 0.0135432f
x_PM_DFFLQNx2_ASAP7_75t_R%MS VSS N_MM11_g N_MM6_d N_MM12_d N_MM7_d N_MM13_d
+ N_MS_3 N_MS_11 N_MS_12 N_MS_13 N_MS_15 N_MS_1 N_MS_17 N_MS_4 N_MS_18 N_MS_14
+ N_MS_16 PM_DFFLQNx2_ASAP7_75t_R%MS
cc_57 N_MS_3 N_CLKN_30 0.000491584f
cc_58 N_MS_3 N_CLKN_10 0.000583016f
cc_59 N_MS_3 N_CLKN_3 0.000123997f
cc_60 N_MS_3 N_MM9_g 0.000162224f
cc_61 N_MS_3 N_CLKN_36 0.000188269f
cc_62 N_MS_11 N_MM12_g 0.00678161f
cc_63 N_MS_12 N_MM12_g 0.00780032f
cc_64 N_MS_13 N_MM12_g 0.00777316f
cc_65 N_MS_15 N_CLKN_10 0.000374991f
cc_66 N_MS_1 N_MM9_g 0.000568369f
cc_67 N_MS_17 N_CLKN_10 0.00153223f
cc_68 N_MS_4 N_MM12_g 0.00231951f
cc_69 N_MS_4 N_CLKN_10 0.00634494f
cc_70 N_MM11_g N_MM9_g 0.0143809f
cc_71 N_MS_3 N_MM12_g 0.0257221f
cc_72 N_MS_13 N_MM10_g 0.000130173f
cc_73 N_MS_13 N_CLKB_19 0.000373469f
cc_74 N_MS_13 N_CLKB_22 0.000205442f
cc_75 N_MS_13 N_CLKB_2 0.000228024f
cc_76 N_MS_17 N_CLKB_19 0.0044299f
cc_77 N_MS_17 N_CLKB_2 0.000385637f
cc_78 N_MS_18 N_CLKB_19 0.000664832f
cc_79 N_MS_14 N_CLKB_22 0.00264321f
cc_80 N_MS_13 N_MM13_g 0.0153919f
x_PM_DFFLQNx2_ASAP7_75t_R%PD2 VSS N_MM10_s N_MM11_d N_PD2_5 N_PD2_1 N_PD2_4
+ PM_DFFLQNx2_ASAP7_75t_R%PD2
cc_81 N_PD2_5 N_CLKN_10 0.00146263f
cc_82 N_PD2_1 N_CLKN_3 0.00052085f
cc_83 N_PD2_1 N_MM9_g 0.00206401f
cc_84 N_PD2_4 N_MM9_g 0.00714445f
cc_85 N_PD2_5 N_MM9_g 0.0240627f
cc_86 N_PD2_4 N_MM10_g 0.0150104f
cc_87 N_PD2_5 N_MM11_g 0.0145937f
cc_88 N_PD2_1 N_MH_16 0.000461869f
cc_89 N_PD2_4 N_MH_3 0.000601241f
cc_90 N_PD2_1 N_MH_20 0.00323624f
x_PM_DFFLQNx2_ASAP7_75t_R%PD5 VSS N_MM17_s N_MM16_d N_PD5_1 N_PD5_4 N_PD5_5
+ PM_DFFLQNx2_ASAP7_75t_R%PD5
cc_91 N_PD5_1 N_MM18_g 0.000859436f
cc_92 N_PD5_4 N_MM18_g 0.00695784f
cc_93 N_PD5_5 N_MM18_g 0.0239997f
cc_94 N_PD5_4 N_MM13_g 0.0153008f
cc_95 N_PD5_1 N_MM19_g 0.000917707f
cc_96 N_PD5_5 N_MM19_g 0.0155867f
cc_97 N_PD5_1 N_SH_14 0.000516396f
cc_98 N_PD5_1 N_SH_16 0.000458254f
cc_99 N_PD5_1 N_SH_17 0.000585951f
cc_100 N_PD5_4 N_SH_5 0.000661838f
cc_101 N_PD5_1 N_SH_25 0.00238444f
x_PM_DFFLQNx2_ASAP7_75t_R%PD1 VSS N_MM5_d N_MM4_s N_PD1_5 N_PD1_4 N_PD1_1
+ PM_DFFLQNx2_ASAP7_75t_R%PD1
cc_102 N_PD1_5 N_CLKN_29 0.000206769f
cc_103 N_PD1_5 N_CLKN_2 0.00209485f
cc_104 N_PD1_5 N_MM1_g 0.0732979f
cc_105 N_PD1_4 N_D_1 0.000671207f
cc_106 N_PD1_4 N_D_4 0.000763833f
cc_107 N_PD1_4 N_MM3_g 0.0361914f
cc_108 N_PD1_5 N_CLKB_18 0.000306126f
cc_109 N_PD1_5 N_CLKB_1 0.000757286f
cc_110 N_PD1_5 N_MM10_g 0.0346069f
cc_111 N_PD1_1 N_MH_4 0.00121056f
cc_112 N_PD1_1 N_MH_10 0.00348783f
x_PM_DFFLQNx2_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_DFFLQNx2_ASAP7_75t_R%noxref_20
cc_113 N_noxref_20_1 N_CLKN_1 0.000129137f
cc_114 N_noxref_20_1 N_MM22_g 0.00352737f
cc_115 N_noxref_20_1 N_CLKB_5 0.000443316f
cc_116 N_noxref_20_1 N_CLKB_13 0.0271608f
x_PM_DFFLQNx2_ASAP7_75t_R%D VSS D N_MM3_g N_D_4 N_D_1 N_D_6 N_D_5
+ PM_DFFLQNx2_ASAP7_75t_R%D
cc_117 N_MM3_g N_CLKN_29 0.000914141f
cc_118 N_D_4 N_CLKN_36 0.000957968f
cc_119 N_D_1 N_CLKN_2 0.00239967f
cc_120 N_D_4 N_CLKN_29 0.00461051f
cc_121 N_MM3_g N_MM1_g 0.00526389f
x_PM_DFFLQNx2_ASAP7_75t_R%SH VSS N_MM14_g N_MM24_g N_MM24@2_g N_MM13_s N_MM18_d
+ N_MM12_s N_MM17_d N_SH_16 N_SH_24 N_SH_26 N_SH_14 N_SH_6 N_SH_19 N_SH_17
+ N_SH_18 N_SH_15 N_SH_5 N_SH_29 N_SH_2 N_SH_23 N_SH_28 N_SH_27 N_SH_21 N_SH_22
+ N_SH_1 N_SH_25 N_SH_20 PM_DFFLQNx2_ASAP7_75t_R%SH
cc_122 N_SH_16 N_CLKN_36 0.00010615f
cc_123 N_SH_24 N_CLKN_10 0.000173239f
cc_124 N_SH_26 N_CLKN_10 0.000204456f
cc_125 N_SH_14 N_MM12_g 0.00677846f
cc_126 N_SH_6 N_CLKN_10 0.000267105f
cc_127 N_SH_19 N_CLKN_5 0.000419009f
cc_128 N_SH_17 N_CLKN_10 0.000429293f
cc_129 N_SH_18 N_CLKN_10 0.00062089f
cc_130 N_SH_15 N_CLKN_5 0.000929177f
cc_131 N_SH_6 N_MM18_g 0.0010039f
cc_132 N_SH_15 N_CLKN_10 0.00226816f
cc_133 N_SH_5 N_MM12_g 0.00951834f
cc_134 N_SH_15 N_MM18_g 0.0162747f
cc_135 N_SH_29 N_CLKB_22 0.000136464f
cc_136 N_SH_6 N_MM13_g 0.000141727f
cc_137 N_SH_19 N_CLKB_19 0.000222283f
cc_138 N_SH_15 N_MM13_g 0.00675261f
cc_139 N_SH_14 N_MM13_g 0.00679213f
cc_140 N_SH_24 N_CLKB_19 0.000311984f
cc_141 N_SH_17 N_CLKB_19 0.00450587f
cc_142 N_SH_17 N_CLKB_2 0.000463902f
cc_143 N_SH_5 N_CLKB_2 0.000532303f
cc_144 N_SH_18 N_CLKB_19 0.000538426f
cc_145 N_SH_26 N_CLKB_19 0.00055759f
cc_146 N_SH_16 N_CLKB_19 0.000565492f
cc_147 N_SH_16 N_CLKB_22 0.00104387f
cc_148 N_SH_5 N_MM13_g 0.0184322f
cc_149 N_SH_18 N_MS_3 0.000109623f
cc_150 N_SH_17 N_MS_3 0.000122722f
cc_151 N_SH_24 N_MS_3 0.000158303f
cc_152 N_SH_15 N_MS_3 0.000437545f
cc_153 N_SH_14 N_MS_3 0.000465191f
cc_154 N_SH_6 N_MS_4 0.000685922f
cc_155 N_SH_24 N_MS_4 0.000297469f
cc_156 N_SH_24 N_MS_17 0.000534102f
cc_157 N_SH_16 N_MS_16 0.000589584f
cc_158 N_SH_15 N_MS_4 0.000599884f
cc_159 N_SH_16 N_MS_18 0.00163826f
cc_160 N_SH_5 N_MS_3 0.00362175f
cc_161 N_SH_16 N_MM19_g 0.000115599f
cc_162 N_SH_18 N_MM19_g 0.000130284f
cc_163 N_SH_2 N_MM19_g 0.000158842f
cc_164 N_SH_23 N_MM19_g 0.000175409f
cc_165 N_SH_28 N_MM19_g 0.000183411f
cc_166 N_SH_27 N_SS_12 0.000219151f
cc_167 N_MM14_g N_SS_10 0.00686383f
cc_168 N_MM14_g N_SS_11 0.00682857f
cc_169 N_SH_21 N_SS_4 0.000249533f
cc_170 N_SH_2 N_SS_15 0.000267699f
cc_171 N_SH_23 N_SS_15 0.00731208f
cc_172 N_SH_22 N_SS_15 0.00182216f
cc_173 N_MM14_g N_SS_3 0.000405f
cc_174 N_MM14_g N_SS_4 0.000527123f
cc_175 N_SH_21 N_SS_14 0.00065136f
cc_176 N_SH_1 N_SS_1 0.00070153f
cc_177 N_SH_25 N_SS_16 0.000793581f
cc_178 N_SH_17 N_SS_1 0.000844674f
cc_179 N_SH_28 N_SS_15 0.000900665f
cc_180 N_SH_20 N_SS_12 0.000954151f
cc_181 N_SH_22 N_SS_13 0.00105941f
cc_182 N_MM14_g N_SS_1 0.00110551f
cc_183 N_SH_1 N_MM19_g 0.00113663f
cc_184 N_SH_28 N_SS_14 0.0012816f
cc_185 N_SH_19 N_SS_12 0.0015353f
cc_186 N_SH_29 N_SS_15 0.00188036f
cc_187 N_SH_17 N_SS_12 0.00474716f
cc_188 N_MM14_g N_MM19_g 0.0293865f
x_PM_DFFLQNx2_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_DFFLQNx2_ASAP7_75t_R%noxref_21
cc_189 N_noxref_21_1 N_CLKN_1 0.000125863f
cc_190 N_noxref_21_1 N_MM22_g 0.00366742f
cc_191 N_noxref_21_1 N_CLKB_6 0.000435904f
cc_192 N_noxref_21_1 N_CLKB_14 0.027101f
cc_193 N_noxref_21_1 N_noxref_20_1 0.00146986f
x_PM_DFFLQNx2_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_DFFLQNx2_ASAP7_75t_R%noxref_22
cc_194 N_noxref_22_1 N_MM3_g 0.00136569f
cc_195 N_noxref_22_1 N_CLKB_13 0.000799075f
cc_196 N_noxref_22_1 N_noxref_20_1 0.00770044f
cc_197 N_noxref_22_1 N_noxref_21_1 0.000471826f
x_PM_DFFLQNx2_ASAP7_75t_R%CLK VSS CLK N_MM20_g N_CLK_8 N_CLK_5 N_CLK_1 N_CLK_6
+ N_CLK_7 N_CLK_4 PM_DFFLQNx2_ASAP7_75t_R%CLK
x_PM_DFFLQNx2_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_DFFLQNx2_ASAP7_75t_R%noxref_23
cc_198 N_noxref_23_1 N_MM3_g 0.0013737f
cc_199 N_noxref_23_1 N_CLKB_14 0.000774644f
cc_200 N_noxref_23_1 N_noxref_20_1 0.000469294f
cc_201 N_noxref_23_1 N_noxref_21_1 0.00769869f
cc_202 N_noxref_23_1 N_noxref_22_1 0.00123377f
x_PM_DFFLQNx2_ASAP7_75t_R%MH VSS N_MM7_g N_MM4_d N_MM9_d N_MM1_d N_MM10_d
+ N_MH_10 N_MH_20 N_MH_3 N_MH_16 N_MH_1 N_MH_17 N_MH_4 N_MH_12 N_MH_14 N_MH_18
+ N_MH_15 N_MH_19 PM_DFFLQNx2_ASAP7_75t_R%MH
cc_203 N_MH_10 N_CLKN_30 0.000373874f
cc_204 N_MH_10 N_MM1_g 0.000402537f
cc_205 N_MH_10 N_CLKN_29 0.000392337f
cc_206 N_MH_20 N_CLKN_30 0.000254895f
cc_207 N_MH_3 N_CLKN_2 0.000280515f
cc_208 N_MH_16 N_CLKN_30 0.00268735f
cc_209 N_MH_1 N_CLKN_10 0.00208847f
cc_210 N_MH_17 N_CLKN_10 0.000621204f
cc_211 N_MH_4 N_MM9_g 0.000631968f
cc_212 N_MH_16 N_CLKN_3 0.000763682f
cc_213 N_MH_12 N_CLKN_2 0.000880938f
cc_214 N_MH_3 N_CLKN_29 0.00133176f
cc_215 N_MH_14 N_CLKN_29 0.00140507f
cc_216 N_MH_14 N_CLKN_36 0.00150368f
cc_217 N_MH_3 N_MM1_g 0.00177621f
cc_218 N_MH_17 N_CLKN_30 0.00361825f
cc_219 N_MM7_g N_CLKN_10 0.00460108f
cc_220 N_MH_12 N_MM1_g 0.0337074f
cc_221 N_MM7_g N_MM12_g 0.0127533f
cc_222 N_MH_10 N_MM9_g 0.0363187f
cc_223 N_MH_10 N_MM13_g 0.00016168f
cc_224 N_MH_10 N_CLKB_18 0.000266136f
cc_225 N_MH_14 N_CLKB_18 0.000329978f
cc_226 N_MH_18 N_CLKB_18 0.00038075f
cc_227 N_MH_12 N_MM10_g 0.0164258f
cc_228 N_MH_3 N_CLKB_1 0.000736382f
cc_229 N_MH_4 N_MM10_g 0.00109557f
cc_230 N_MH_15 N_CLKB_18 0.00111855f
cc_231 N_MH_3 N_MM10_g 0.00117424f
cc_232 N_MH_17 N_CLKB_22 0.00124947f
cc_233 N_MH_16 N_CLKB_18 0.00135198f
cc_234 N_MH_12 N_CLKB_1 0.0018255f
cc_235 N_MH_16 N_CLKB_22 0.00226638f
cc_236 N_MH_19 N_CLKB_18 0.00273185f
cc_237 N_MH_10 N_MM10_g 0.0530885f
cc_238 N_MH_4 N_MS_1 0.000401853f
cc_239 N_MH_17 N_MS_18 0.000564126f
cc_240 N_MH_17 N_MS_1 0.000830281f
cc_241 N_MH_1 N_MS_14 0.000836487f
cc_242 N_MH_17 N_MS_17 0.000959232f
cc_243 N_MM7_g N_MS_3 0.000974987f
cc_244 N_MH_1 N_MM11_g 0.00106092f
cc_245 N_MM7_g N_MS_1 0.00116111f
cc_246 N_MH_15 N_MS_14 0.0012402f
cc_247 N_MM7_g N_MS_12 0.0063972f
cc_248 N_MM7_g N_MS_11 0.00641046f
cc_249 N_MH_17 N_MS_14 0.00719325f
cc_250 N_MM7_g N_MM11_g 0.0293111f
x_PM_DFFLQNx2_ASAP7_75t_R%CLKN VSS N_MM22_g N_MM1_g N_MM9_g N_MM12_g N_MM18_g
+ N_MM20_d N_MM21_d N_CLKN_28 N_CLKN_35 N_CLKN_32 N_CLKN_9 N_CLKN_34 N_CLKN_8
+ N_CLKN_21 N_CLKN_22 N_CLKN_26 N_CLKN_25 N_CLKN_1 N_CLKN_27 N_CLKN_36
+ N_CLKN_23 N_CLKN_29 N_CLKN_2 N_CLKN_5 N_CLKN_30 N_CLKN_3 N_CLKN_10 N_CLKN_31
+ N_CLKN_33 N_CLKN_24 PM_DFFLQNx2_ASAP7_75t_R%CLKN
cc_251 N_CLKN_28 N_MM20_g 8.64818e-20
cc_252 N_CLKN_35 N_MM20_g 8.69563e-20
cc_253 N_CLKN_32 N_MM20_g 0.000192798f
cc_254 N_CLKN_9 N_MM20_g 0.00109915f
cc_255 N_CLKN_34 N_MM20_g 0.000233607f
cc_256 N_CLKN_8 N_MM20_g 0.00117509f
cc_257 N_CLKN_21 N_MM20_g 0.0112203f
cc_258 N_CLKN_22 N_MM20_g 0.0113257f
cc_259 N_CLKN_26 N_CLK_8 0.000734123f
cc_260 N_CLKN_25 N_CLK_5 0.000758513f
cc_261 N_CLKN_1 N_CLK_8 0.000777867f
cc_262 N_CLKN_27 N_CLK_1 0.000922771f
cc_263 N_CLKN_26 N_CLK_6 0.00131231f
cc_264 N_CLKN_27 N_CLK_7 0.0013657f
cc_265 N_CLKN_36 N_CLK_8 0.0016944f
cc_266 N_CLKN_23 N_CLK_4 0.00176132f
cc_267 N_CLKN_27 N_CLK_4 0.00214909f
cc_268 N_CLKN_34 N_CLK_8 0.00227131f
cc_269 N_CLKN_25 N_CLK_7 0.00227493f
cc_270 N_CLKN_1 N_CLK_1 0.00232584f
cc_271 N_CLKN_27 N_CLK_8 0.00241801f
cc_272 N_CLKN_32 N_CLK_8 0.00279116f
cc_273 N_MM22_g N_MM20_g 0.0351395f
x_PM_DFFLQNx2_ASAP7_75t_R%CLKB VSS N_MM10_g N_MM13_g N_MM23_d N_MM22_d
+ N_CLKB_17 N_CLKB_6 N_CLKB_5 N_CLKB_16 N_CLKB_15 N_CLKB_13 N_CLKB_21 N_CLKB_22
+ N_CLKB_14 N_CLKB_19 N_CLKB_18 N_CLKB_2 N_CLKB_1 N_CLKB_20
+ PM_DFFLQNx2_ASAP7_75t_R%CLKB
cc_274 N_CLKB_17 N_CLK_5 9.42661e-20
cc_275 N_CLKB_6 N_CLK_5 0.000321239f
cc_276 N_CLKB_5 N_CLK_5 0.000406233f
cc_277 N_CLKB_16 N_CLK_5 0.000213606f
cc_278 N_CLKB_16 N_CLK_6 0.000974336f
cc_279 N_CLKB_15 N_CLK_5 0.00220356f
cc_280 N_CLKB_13 N_CLKN_26 3.22363e-20
cc_281 N_CLKB_13 N_CLKN_23 6.36253e-20
cc_282 N_MM13_g N_CLKN_5 0.000222584f
cc_283 N_CLKB_21 N_CLKN_34 0.000231065f
cc_284 N_CLKB_6 N_CLKN_34 0.000271072f
cc_285 N_CLKB_22 N_CLKN_30 0.000665549f
cc_286 N_CLKB_6 N_CLKN_1 0.000308943f
cc_287 N_CLKB_14 N_MM22_g 0.0112471f
cc_288 N_CLKB_16 N_CLKN_34 0.00508495f
cc_289 N_CLKB_22 N_CLKN_29 0.000355479f
cc_290 N_CLKB_15 N_CLKN_35 0.000457217f
cc_291 N_MM10_g N_CLKN_3 0.000540881f
cc_292 N_CLKB_19 N_CLKN_10 0.000573176f
cc_293 N_CLKB_18 N_CLKN_36 0.000611247f
cc_294 N_CLKB_14 N_CLKN_1 0.000622622f
cc_295 N_CLKB_6 N_CLKN_27 0.000664076f
cc_296 N_CLKB_2 N_CLKN_10 0.00285577f
cc_297 N_CLKB_17 N_CLKN_36 0.000735061f
cc_298 N_CLKB_5 N_MM22_g 0.000758246f
cc_299 N_CLKB_1 N_CLKN_2 0.00227225f
cc_300 N_CLKB_17 N_CLKN_28 0.000987161f
cc_301 N_CLKB_6 N_MM22_g 0.00107449f
cc_302 N_MM10_g N_MM1_g 0.00162813f
cc_303 N_CLKB_18 N_CLKN_29 0.00310318f
cc_304 N_CLKB_17 N_CLKN_35 0.00376577f
cc_305 N_MM13_g N_CLKN_10 0.00430634f
cc_306 N_MM13_g N_MM12_g 0.00567108f
cc_307 N_MM10_g N_MM9_g 0.00910719f
cc_308 N_MM13_g N_MM18_g 0.0184479f
cc_309 N_CLKB_22 N_CLKN_36 0.0282547f
cc_310 N_CLKB_13 N_MM22_g 0.03884f
cc_311 N_CLKB_18 N_D_4 0.000146015f
cc_312 N_CLKB_21 N_D_6 0.000777105f
cc_313 N_CLKB_20 N_D_5 0.00096655f
cc_314 N_CLKB_22 N_D_4 0.00108401f
cc_315 N_CLKB_17 N_D_4 0.0083886f
*END of DFFLQNx2_ASAP7_75t_R.pxi
.ENDS
** Design:	DFFLQNx3_ASAP7_75t_R
* Created:	"Fri Aug 17 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "DFFLQNx3_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "DFFLQNx3_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_DFFLQNx3_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.0418508f
.ends

.subckt PM_DFFLQNx3_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.0418132f
.ends

.subckt PM_DFFLQNx3_ASAP7_75t_R%PD4 VSS 2 4 1
c1 1 VSS 0.000948557f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.2295 $X2=0.7605 $Y2=0.2295
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.2295 $X2=0.7435 $Y2=0.2295
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7435 $Y=0.2295 $X2=0.7605 $Y2=0.2295
.ends

.subckt PM_DFFLQNx3_ASAP7_75t_R%PD3 VSS 2 4 1
c1 1 VSS 0.000983844f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0405 $X2=0.4905 $Y2=0.0405
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0405 $X2=0.4735 $Y2=0.0405
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4735 $Y=0.0405 $X2=0.4905 $Y2=0.0405
.ends

.subckt PM_DFFLQNx3_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.00418573f
.ends

.subckt PM_DFFLQNx3_ASAP7_75t_R%PU1 VSS 2 4 1
c1 1 VSS 0.000973869f
r1 4 3 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3365 $Y2=0.2025
r2 2 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3195 $Y2=0.2025
r3 1 3 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3195 $Y=0.2025 $X2=0.3365 $Y2=0.2025
.ends

.subckt PM_DFFLQNx3_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.00417063f
.ends

.subckt PM_DFFLQNx3_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.00470193f
.ends

.subckt PM_DFFLQNx3_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.00478217f
.ends

.subckt PM_DFFLQNx3_ASAP7_75t_R%PD2 VSS 7 12 5 1 4
c1 1 VSS 0.00727636f
c2 4 VSS 0.00188706f
c3 5 VSS 0.00233436f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4880 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r3 9 5 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.4605
+ $Y=0.2295 $X2=0.4860 $Y2=0.2295
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.4455
+ $Y=0.2295 $X2=0.4605 $Y2=0.2295
r5 1 8 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4320
+ $Y=0.2295 $X2=0.4455 $Y2=0.2295
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2295 $X2=0.4300 $Y2=0.2295
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2295 $X2=0.4175 $Y2=0.2295
.ends

.subckt PM_DFFLQNx3_ASAP7_75t_R%PD1 VSS 7 10 5 4 1
c1 1 VSS 0.0097274f
c2 4 VSS 0.00316998f
c3 5 VSS 0.00186047f
r1 10 9 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r2 8 9 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r3 5 8 0.123457 $w=8.1e-08 $l=1e-08 $layer=N_src_drn $thickness=1e-09 $X=0.3780
+ $Y=0.0675 $X2=0.3880 $Y2=0.0675
r4 4 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3220 $Y2=0.0675
r5 7 4 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r6 1 5 1e-05
.ends

.subckt PM_DFFLQNx3_ASAP7_75t_R%D VSS 9 3 4 1 6 5
c1 1 VSS 0.00681633f
c2 3 VSS 0.0834273f
c3 4 VSS 0.00585921f
c4 5 VSS 0.00683405f
c5 6 VSS 0.00763269f
r1 6 13 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.2340 $X2=0.2970 $Y2=0.2140
r2 5 8 5.17411 $w=1.46514e-08 $l=2.72e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0360 $X2=0.2970 $Y2=0.0632
r3 12 13 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1735 $X2=0.2970 $Y2=0.2140
r4 11 12 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1735
r5 9 10 2.85657 $w=1.3e-08 $l=1.22e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0820 $X2=0.2970 $Y2=0.0942
r6 9 8 4.37231 $w=1.3e-08 $l=1.88e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0820 $X2=0.2970 $Y2=0.0632
r7 4 10 5.07188 $w=1.3e-08 $l=2.18e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1160 $X2=0.2970 $Y2=0.0942
r8 4 11 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1160 $X2=0.2970 $Y2=0.1350
r9 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r10 1 11 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_DFFLQNx3_ASAP7_75t_R%CLK VSS 11 3 8 5 1 6 7 4
c1 1 VSS 0.00261608f
c2 3 VSS 0.0598018f
c3 4 VSS 0.001052f
c4 5 VSS 0.0041429f
c5 6 VSS 0.00373722f
c6 7 VSS 0.00235054f
c7 8 VSS 0.00198788f
r1 6 17 3.22357 $w=2.26279e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.2125 $X2=0.1080 $Y2=0.1820
r2 5 15 3.22357 $w=2.26279e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0575 $X2=0.1080 $Y2=0.0880
r3 16 17 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.1820 $X2=0.1080 $Y2=0.1820
r4 8 13 2.6406 $w=2.38947e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1820 $X2=0.0810 $Y2=0.1540
r5 8 16 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1820 $X2=0.0945 $Y2=0.1820
r6 14 15 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.0880 $X2=0.1080 $Y2=0.0880
r7 7 10 1.76614 $w=2.65738e-08 $l=2.42e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0880 $X2=0.0810 $Y2=0.1122
r8 7 14 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0880 $X2=0.0945 $Y2=0.0880
r9 11 12 0.874462 $w=1.3e-08 $l=3.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1227
r10 11 10 1.57403 $w=1.3e-08 $l=6.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1122
r11 4 12 2.85657 $w=1.3e-08 $l=1.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1227
r12 4 13 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1540
r13 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r14 1 4 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_DFFLQNx3_ASAP7_75t_R%MH VSS 9 47 51 57 61 10 20 3 16 1 17 4 12 14 18
+ 15 19
c1 1 VSS 0.000275646f
c2 3 VSS 0.00624319f
c3 4 VSS 0.00540796f
c4 9 VSS 0.0363983f
c5 10 VSS 0.00227021f
c6 11 VSS 8.98741e-20
c7 12 VSS 0.00278014f
c8 13 VSS 6.87463e-20
c9 14 VSS 0.00852088f
c10 15 VSS 0.00125663f
c11 16 VSS 0.000667671f
c12 17 VSS 0.000549286f
c13 18 VSS 0.00649583f
c14 19 VSS 1.21134e-20
c15 20 VSS 0.00228279f
r1 61 60 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r2 59 60 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r3 3 59 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3760 $Y=0.2295 $X2=0.3880 $Y2=0.2295
r4 13 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2295 $X2=0.3760 $Y2=0.2295
r5 55 56 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r6 57 55 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.1890 $X2=0.3635 $Y2=0.1890
r7 12 56 0.185185 $w=5.4e-08 $l=1e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r8 12 3 0.518519 $w=3.9e-08 $l=4.05494e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.1890 $X2=0.3760 $Y2=0.2295
r9 3 44 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2295
+ $X2=0.3780 $Y2=0.2340
r10 51 50 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r11 49 50 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4420 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r12 4 49 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4300 $Y=0.0405 $X2=0.4420 $Y2=0.0405
r13 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0405 $X2=0.4300 $Y2=0.0405
r14 10 4 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0810 $X2=0.4300 $Y2=0.0810
r15 47 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0810 $X2=0.4175 $Y2=0.0810
r16 44 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r17 42 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r18 41 42 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4160
+ $Y=0.2340 $X2=0.4050 $Y2=0.2340
r19 14 20 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4340
+ $Y=0.2340 $X2=0.4590 $Y2=0.2340
r20 14 41 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4340
+ $Y=0.2340 $X2=0.4160 $Y2=0.2340
r21 4 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0405
+ $X2=0.4320 $Y2=0.0360
r22 20 34 3.01468 $w=1.741e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4590 $Y2=0.2140
r23 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4455 $Y2=0.0360
r24 18 31 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4590 $Y2=0.0630
r25 18 37 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4455 $Y2=0.0360
r26 33 34 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1850 $X2=0.4590 $Y2=0.2140
r27 32 33 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1660 $X2=0.4590 $Y2=0.1850
r28 16 19 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1525 $X2=0.4590 $Y2=0.1310
r29 16 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1525 $X2=0.4590 $Y2=0.1660
r30 30 31 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0900 $X2=0.4590 $Y2=0.0630
r31 29 30 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1025 $X2=0.4590 $Y2=0.0900
r32 15 19 2.78392 $w=1.56471e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1140 $X2=0.4590 $Y2=0.1310
r33 15 29 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1140 $X2=0.4590 $Y2=0.1025
r34 19 27 4.18306 $w=1.49565e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1310 $X2=0.4820 $Y2=0.1310
r35 26 27 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5000
+ $Y=0.1310 $X2=0.4820 $Y2=0.1310
r36 25 26 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1310 $X2=0.5000 $Y2=0.1310
r37 17 24 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1310 $X2=0.5670 $Y2=0.1310
r38 17 25 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1310 $X2=0.5130 $Y2=0.1310
r39 23 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1330
+ $X2=0.5670 $Y2=0.1310
r40 1 22 1.47681 $w=1.53e-08 $l=9e-09 $layer=LIG $thickness=4.8e-08 $X=0.5670
+ $Y=0.1215 $X2=0.5670 $Y2=0.1305
r41 22 23 5.31651 $w=1.53e-08 $l=2.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.5670 $Y=0.1305 $X2=0.5670 $Y2=0.1330
r42 9 22 0.314665 $w=2.27e-07 $l=4.5e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5670 $Y=0.1350 $X2=0.5670 $Y2=0.1305
r43 3 12 1e-05
.ends

.subckt PM_DFFLQNx3_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.0042337f
.ends

.subckt PM_DFFLQNx3_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.00431915f
.ends

.subckt PM_DFFLQNx3_ASAP7_75t_R%SS VSS 9 31 40 12 10 11 4 15 3 14 1 16 13
c1 1 VSS 0.00107305f
c2 3 VSS 0.00625569f
c3 4 VSS 0.00661472f
c4 9 VSS 0.0384302f
c5 10 VSS 0.00321334f
c6 11 VSS 0.00319596f
c7 12 VSS 0.00183358f
c8 13 VSS 0.0137221f
c9 14 VSS 0.00921325f
c10 15 VSS 0.00698424f
c11 16 VSS 0.00323748f
c12 17 VSS 0.00348834f
c13 18 VSS 0.00345666f
r1 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.2295 $X2=0.8620 $Y2=0.2295
r2 40 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.2295 $X2=0.8495 $Y2=0.2295
r3 4 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.2295
+ $X2=0.8640 $Y2=0.2340
r4 37 38 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.2340 $X2=0.8865 $Y2=0.2340
r5 14 18 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9180 $Y=0.2340 $X2=0.9450 $Y2=0.2340
r6 14 38 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.2340 $X2=0.8865 $Y2=0.2340
r7 18 35 6.74572 $w=1.545e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.2340 $X2=0.9450 $Y2=0.1980
r8 34 35 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1690 $X2=0.9450 $Y2=0.1980
r9 33 34 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1420 $X2=0.9450 $Y2=0.1690
r10 32 33 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1035 $X2=0.9450 $Y2=0.1420
r11 15 17 5.69636 $w=1.58e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.0675 $X2=0.9450 $Y2=0.0360
r12 15 32 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.0675 $X2=0.9450 $Y2=0.1035
r13 10 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.0405 $X2=0.8620 $Y2=0.0405
r14 31 10 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.0405 $X2=0.8495 $Y2=0.0405
r15 17 29 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.0360 $X2=0.9180 $Y2=0.0360
r16 3 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.0405
+ $X2=0.8640 $Y2=0.0360
r17 28 29 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.0360 $X2=0.9180 $Y2=0.0360
r18 27 28 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.0360 $X2=0.8910 $Y2=0.0360
r19 26 27 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.0360 $X2=0.8640 $Y2=0.0360
r20 13 16 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.0360 $X2=0.7830 $Y2=0.0360
r21 13 26 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0360 $X2=0.8370 $Y2=0.0360
r22 12 23 8.04505 $w=1.3e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.0705 $X2=0.7830 $Y2=0.1050
r23 12 16 6.39593 $w=1.55565e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7830 $Y=0.0705 $X2=0.7830 $Y2=0.0360
r24 1 20 2.36633 $w=2.3e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.7830
+ $Y=0.1055 $X2=0.7830 $Y2=0.1055
r25 1 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7830 $Y=0.1055
+ $X2=0.7830 $Y2=0.1050
r26 9 20 0.314665 $w=2.27e-07 $l=2.95e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.7830 $Y=0.1350 $X2=0.7830 $Y2=0.1055
.ends

.subckt PM_DFFLQNx3_ASAP7_75t_R%PD5 VSS 7 12 1 4 5
c1 1 VSS 0.00746579f
c2 4 VSS 0.00187606f
c3 5 VSS 0.00237762f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.0405 $X2=0.7705 $Y2=0.0405
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7580 $Y=0.0405 $X2=0.7705 $Y2=0.0405
r3 9 5 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.7425
+ $Y=0.0405 $X2=0.7560 $Y2=0.0405
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.7275
+ $Y=0.0405 $X2=0.7425 $Y2=0.0405
r5 1 8 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.7020
+ $Y=0.0405 $X2=0.7275 $Y2=0.0405
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.0405 $X2=0.7000 $Y2=0.0405
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.0405 $X2=0.6875 $Y2=0.0405
.ends

.subckt PM_DFFLQNx3_ASAP7_75t_R%noxref_28 VSS 1
c1 1 VSS 0.00558846f
.ends

.subckt PM_DFFLQNx3_ASAP7_75t_R%noxref_26 VSS 1
c1 1 VSS 0.0414822f
.ends

.subckt PM_DFFLQNx3_ASAP7_75t_R%noxref_27 VSS 1
c1 1 VSS 0.0414795f
.ends

.subckt PM_DFFLQNx3_ASAP7_75t_R%QN VSS 32 24 25 36 43 44 46 13 19 18 15 3 4 1 2
+ 16 14
c1 1 VSS 0.0103125f
c2 2 VSS 0.0112258f
c3 3 VSS 0.00800469f
c4 4 VSS 0.00781134f
c5 13 VSS 0.00456492f
c6 14 VSS 0.00344614f
c7 15 VSS 0.00454848f
c8 16 VSS 0.00344414f
c9 17 VSS 0.0146027f
c10 18 VSS 0.0145552f
c11 19 VSS 0.00374519f
c12 20 VSS 0.00270931f
c13 21 VSS 0.00271104f
r1 16 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.1195 $Y=0.2025 $X2=1.1320 $Y2=0.2025
r2 46 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.1170 $Y=0.2025 $X2=1.1195 $Y2=0.2025
r3 44 42 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0430 $Y=0.2025 $X2=1.0405 $Y2=0.2025
r4 2 42 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0260 $Y=0.2025 $X2=1.0405 $Y2=0.2025
r5 15 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0115 $Y=0.2025 $X2=1.0260 $Y2=0.2025
r6 43 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0090 $Y=0.2025 $X2=1.0115 $Y2=0.2025
r7 4 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.1340 $Y=0.2025
+ $X2=1.1340 $Y2=0.2340
r8 2 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0260 $Y=0.2025
+ $X2=1.0260 $Y2=0.2340
r9 39 40 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.1340
+ $Y=0.2340 $X2=1.1480 $Y2=0.2340
r10 38 39 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.0800
+ $Y=0.2340 $X2=1.1340 $Y2=0.2340
r11 37 38 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.2340 $X2=1.0800 $Y2=0.2340
r12 18 37 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.0145
+ $Y=0.2340 $X2=1.0260 $Y2=0.2340
r13 21 34 7.2121 $w=1.53211e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1620 $Y=0.2340 $X2=1.1620 $Y2=0.1960
r14 21 40 1.61554 $w=1.62143e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1620 $Y=0.2340 $X2=1.1480 $Y2=0.2340
r15 14 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.1195 $Y=0.0675 $X2=1.1320 $Y2=0.0675
r16 36 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.1170 $Y=0.0675 $X2=1.1195 $Y2=0.0675
r17 33 34 11.1348 $w=1.3e-08 $l=4.78e-08 $layer=M1 $thickness=3.6e-08 $X=1.1620
+ $Y=0.1482 $X2=1.1620 $Y2=0.1960
r18 32 33 4.4889 $w=1.3e-08 $l=1.92e-08 $layer=M1 $thickness=3.6e-08 $X=1.1620
+ $Y=0.1290 $X2=1.1620 $Y2=0.1482
r19 32 31 4.6055 $w=1.3e-08 $l=1.98e-08 $layer=M1 $thickness=3.6e-08 $X=1.1620
+ $Y=0.1290 $X2=1.1620 $Y2=0.1092
r20 19 20 5.69636 $w=1.58e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1620 $Y=0.0675 $X2=1.1620 $Y2=0.0360
r21 19 31 9.73567 $w=1.3e-08 $l=4.17e-08 $layer=M1 $thickness=3.6e-08 $X=1.1620
+ $Y=0.0675 $X2=1.1620 $Y2=0.1092
r22 3 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.1340 $Y=0.0675
+ $X2=1.1340 $Y2=0.0360
r23 20 30 1.61554 $w=1.62143e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1620 $Y=0.0360 $X2=1.1480 $Y2=0.0360
r24 29 30 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.1340
+ $Y=0.0360 $X2=1.1480 $Y2=0.0360
r25 28 29 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.0800
+ $Y=0.0360 $X2=1.1340 $Y2=0.0360
r26 27 28 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.0360 $X2=1.0800 $Y2=0.0360
r27 26 27 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.0145
+ $Y=0.0360 $X2=1.0260 $Y2=0.0360
r28 17 26 0.699569 $w=1.3e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=1.0115
+ $Y=0.0360 $X2=1.0145 $Y2=0.0360
r29 1 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0260 $Y=0.0675
+ $X2=1.0260 $Y2=0.0360
r30 25 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.0430 $Y=0.0675 $X2=1.0405 $Y2=0.0675
r31 1 23 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.0260 $Y=0.0675 $X2=1.0405 $Y2=0.0675
r32 13 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.0115 $Y=0.0675 $X2=1.0260 $Y2=0.0675
r33 24 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.0090 $Y=0.0675 $X2=1.0115 $Y2=0.0675
.ends

.subckt PM_DFFLQNx3_ASAP7_75t_R%CLKN VSS 16 17 18 19 20 99 101 28 35 32 9 34 8
+ 21 22 26 25 1 27 36 23 29 2 5 30 3 10 31 33 24
c1 1 VSS 0.0014837f
c2 2 VSS 0.000298835f
c3 3 VSS 7.26317e-20
c4 4 VSS 1e-36
c5 5 VSS 0.000412935f
c6 8 VSS 0.00771637f
c7 9 VSS 0.00772058f
c8 10 VSS 0.00355123f
c9 16 VSS 0.0590851f
c10 17 VSS 0.00560956f
c11 18 VSS 0.005115f
c12 19 VSS 0.0043807f
c13 20 VSS 0.00518077f
c14 21 VSS 0.00657473f
c15 22 VSS 0.00652508f
c16 23 VSS 0.00802558f
c17 24 VSS 0.00181301f
c18 25 VSS 0.00454572f
c19 26 VSS 0.00375681f
c20 27 VSS 0.000659046f
c21 28 VSS 0.000261303f
c22 29 VSS 0.000827386f
c23 30 VSS 0.00146415f
c24 31 VSS 0.00383798f
c25 32 VSS 0.00190812f
c26 33 VSS 0.00393829f
c27 34 VSS 0.000841979f
c28 35 VSS 0.000478248f
c29 36 VSS 0.0227838f
r1 101 100 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r2 22 100 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r3 99 98 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r4 21 98 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r5 9 96 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0550 $Y2=0.2340
r6 8 93 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0550 $Y2=0.0360
r7 95 96 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.2340 $X2=0.0550 $Y2=0.2340
r8 26 95 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0460 $Y2=0.2340
r9 26 33 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0180 $Y2=0.2340
r10 92 93 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.0360 $X2=0.0550 $Y2=0.0360
r11 25 92 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0460 $Y2=0.0360
r12 25 31 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0180 $Y2=0.0360
r13 5 91 2.78395 $w=2.4e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08 $X=0.7290
+ $Y=0.1780 $X2=0.7250 $Y2=0.1780
r14 20 5 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.7290 $Y=0.1350 $X2=0.7290 $Y2=0.1780
r15 4 84 10.3807 $w=2.30357e-08 $l=0 $layer=LISD $thickness=3.675e-08 $X=0.6210
+ $Y=0.1780 $X2=0.6210 $Y2=0.1780
r16 19 4 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.6210 $Y=0.1350 $X2=0.6210 $Y2=0.1780
r17 3 77 2.78395 $w=2.4e-08 $l=5e-09 $layer=LIG $thickness=4.8e-08 $X=0.4590
+ $Y=0.1780 $X2=0.4640 $Y2=0.1780
r18 18 3 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4590 $Y2=0.1780
r19 33 72 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.2340 $X2=0.0180 $Y2=0.2125
r20 31 71 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.0360 $X2=0.0180 $Y2=0.0575
r21 90 91 4.8113 $w=2.22e-08 $l=1.5e-09 $layer=LISD $thickness=2.7e-08
+ $X=0.7235 $Y=0.1780 $X2=0.7250 $Y2=0.1780
r22 89 90 10.8887 $w=2.22e-08 $l=2.15e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7020 $Y=0.1780 $X2=0.7235 $Y2=0.1780
r23 88 89 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6885 $Y=0.1780 $X2=0.7020 $Y2=0.1780
r24 87 88 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6750 $Y=0.1780 $X2=0.6885 $Y2=0.1780
r25 86 87 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6615 $Y=0.1780 $X2=0.6750 $Y2=0.1780
r26 85 86 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6480 $Y=0.1780 $X2=0.6615 $Y2=0.1780
r27 84 85 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6210 $Y=0.1780 $X2=0.6480 $Y2=0.1780
r28 83 84 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5940 $Y=0.1780 $X2=0.6210 $Y2=0.1780
r29 82 83 7.09034 $w=2.22e-08 $l=1.4e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5800 $Y=0.1780 $X2=0.5940 $Y2=0.1780
r30 81 82 6.58388 $w=2.22e-08 $l=1.3e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5670 $Y=0.1780 $X2=0.5800 $Y2=0.1780
r31 80 81 6.58388 $w=2.22e-08 $l=1.3e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5540 $Y=0.1780 $X2=0.5670 $Y2=0.1780
r32 79 80 7.09034 $w=2.22e-08 $l=1.4e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5400 $Y=0.1780 $X2=0.5540 $Y2=0.1780
r33 78 79 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5265 $Y=0.1780 $X2=0.5400 $Y2=0.1780
r34 76 77 10.3823 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4775 $Y=0.1780 $X2=0.4640 $Y2=0.1780
r35 75 76 11.142 $w=2.22e-08 $l=2.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4995 $Y=0.1780 $X2=0.4775 $Y2=0.1780
r36 74 78 1.51936 $w=2.22e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.5235
+ $Y=0.1780 $X2=0.5265 $Y2=0.1780
r37 73 74 5.31775 $w=2.22e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5130 $Y=0.1780 $X2=0.5235 $Y2=0.1780
r38 10 73 5.31775 $w=2.22e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5025 $Y=0.1780 $X2=0.5130 $Y2=0.1780
r39 10 75 1.51936 $w=2.22e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.5025
+ $Y=0.1780 $X2=0.4995 $Y2=0.1780
r40 2 65 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
r41 17 2 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r42 24 32 0.998523 $w=1.74118e-08 $l=1.01119e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1990 $X2=0.0165 $Y2=0.1890
r43 24 72 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1990 $X2=0.0180 $Y2=0.2125
r44 70 71 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0880 $X2=0.0180 $Y2=0.0575
r45 69 70 10.9599 $w=1.3e-08 $l=4.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1350 $X2=0.0180 $Y2=0.0880
r46 23 32 2.63085 $w=1.54194e-08 $l=1.7066e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1720 $X2=0.0165 $Y2=0.1890
r47 23 69 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1720 $X2=0.0180 $Y2=0.1350
r48 67 73 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5130 $Y=0.1845
+ $X2=0.5130 $Y2=0.1780
r49 30 67 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1680 $X2=0.5130 $Y2=0.1845
r50 65 66 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1555
r51 29 63 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1735 $X2=0.3510 $Y2=0.1890
r52 29 66 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1735 $X2=0.3510 $Y2=0.1555
r53 60 61 1.90199 $w=1.38333e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.0255 $Y=0.1890 $X2=0.0345 $Y2=0.1890
r54 32 60 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0165
+ $Y=0.1890 $X2=0.0255 $Y2=0.1890
r55 58 67 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.5130 $Y=0.1890
+ $X2=0.5130 $Y2=0.1845
r56 57 58 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.4320
+ $Y=0.1890 $X2=0.5130 $Y2=0.1890
r57 56 57 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1890 $X2=0.4320 $Y2=0.1890
r58 56 63 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.3510 $Y=0.1890
+ $X2=0.3510 $Y2=0.1890
r59 55 56 15.2739 $w=1.3e-08 $l=6.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.2855
+ $Y=0.1890 $X2=0.3510 $Y2=0.1890
r60 54 55 20.2875 $w=1.3e-08 $l=8.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.1985
+ $Y=0.1890 $X2=0.2855 $Y2=0.1890
r61 53 54 9.211 $w=1.3e-08 $l=3.95e-08 $layer=M2 $thickness=3.6e-08 $X=0.1590
+ $Y=0.1890 $X2=0.1985 $Y2=0.1890
r62 52 53 14.691 $w=1.3e-08 $l=6.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.0960
+ $Y=0.1890 $X2=0.1590 $Y2=0.1890
r63 51 52 14.691 $w=1.3e-08 $l=6.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.0330
+ $Y=0.1890 $X2=0.0960 $Y2=0.1890
r64 51 61 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.0330 $Y=0.1890
+ $X2=0.0345 $Y2=0.1890
r65 36 51 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.0215
+ $Y=0.1890 $X2=0.0330 $Y2=0.1890
r66 48 49 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1590
+ $Y=0.1890 $X2=0.1740 $Y2=0.1890
r67 48 53 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1590 $Y=0.1890
+ $X2=0.1590 $Y2=0.1890
r68 34 46 2.78392 $w=1.56471e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1890 $X2=0.1890 $Y2=0.1720
r69 34 49 2.31754 $w=1.6e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1890 $X2=0.1740 $Y2=0.1890
r70 28 35 2.78149 $w=1.76421e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1540 $X2=0.1890 $Y2=0.1350
r71 28 46 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1540 $X2=0.1890 $Y2=0.1720
r72 35 45 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1640 $Y2=0.1350
r73 44 45 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.1465
+ $Y=0.1350 $X2=0.1640 $Y2=0.1350
r74 43 44 0.46638 $w=1.3e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.1445
+ $Y=0.1350 $X2=0.1465 $Y2=0.1350
r75 42 43 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1445 $Y2=0.1350
r76 27 42 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1235
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r77 16 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r78 1 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
r79 9 22 1e-05
r80 8 21 1e-05
.ends

.subckt PM_DFFLQNx3_ASAP7_75t_R%MS VSS 10 39 42 47 49 3 11 12 13 15 1 17 4 18
+ 14 16
c1 1 VSS 0.00219677f
c2 3 VSS 0.0053734f
c3 4 VSS 0.00934756f
c4 10 VSS 0.0375014f
c5 11 VSS 0.0028652f
c6 12 VSS 0.00269664f
c7 13 VSS 0.00225966f
c8 14 VSS 0.00187004f
c9 15 VSS 0.00403627f
c10 16 VSS 0.00299125f
c11 17 VSS 0.00103806f
c12 18 VSS 0.000436471f
c13 19 VSS 0.00295242f
r1 49 48 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.2295 $X2=0.6625 $Y2=0.2295
r2 13 48 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6500 $Y=0.2295 $X2=0.6625 $Y2=0.2295
r3 12 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2295 $X2=0.5920 $Y2=0.2295
r4 47 12 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.2295 $X2=0.5795 $Y2=0.2295
r5 44 13 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6210 $Y=0.2295 $X2=0.6480 $Y2=0.2295
r6 4 44 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08 $X=0.5940
+ $Y=0.2295 $X2=0.6210 $Y2=0.2295
r7 4 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2295
+ $X2=0.5965 $Y2=0.2340
r8 15 19 4.06404 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5965 $Y=0.2340 $X2=0.6210 $Y2=0.2340
r9 42 41 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.0405 $X2=0.6085 $Y2=0.0405
r10 40 41 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6040 $Y=0.0405 $X2=0.6085 $Y2=0.0405
r11 3 40 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5920 $Y=0.0405 $X2=0.6040 $Y2=0.0405
r12 11 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.0405 $X2=0.5920 $Y2=0.0405
r13 39 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0405 $X2=0.5795 $Y2=0.0405
r14 19 35 3.01468 $w=1.741e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.2340 $X2=0.6210 $Y2=0.2140
r15 3 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0405
+ $X2=0.5940 $Y2=0.0540
r16 34 35 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1850 $X2=0.6210 $Y2=0.2140
r17 33 34 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1660 $X2=0.6210 $Y2=0.1850
r18 32 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1525 $X2=0.6210 $Y2=0.1660
r19 31 32 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1310 $X2=0.6210 $Y2=0.1525
r20 17 28 3.60008 $w=1.51951e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.1105 $X2=0.6210 $Y2=0.0900
r21 17 31 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1105 $X2=0.6210 $Y2=0.1310
r22 16 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0540 $X2=0.5940 $Y2=0.0720
r23 27 28 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6075 $Y=0.0900 $X2=0.6210 $Y2=0.0900
r24 18 26 1.38478 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5940 $Y=0.0900 $X2=0.5830 $Y2=0.0900
r25 18 27 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5940 $Y=0.0900 $X2=0.6075 $Y2=0.0900
r26 18 29 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0900 $X2=0.5940 $Y2=0.0720
r27 25 26 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5515
+ $Y=0.0900 $X2=0.5830 $Y2=0.0900
r28 24 25 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0900 $X2=0.5515 $Y2=0.0900
r29 14 24 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5000
+ $Y=0.0900 $X2=0.5130 $Y2=0.0900
r30 1 21 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.5130
+ $Y=0.0900 $X2=0.5130 $Y2=0.0900
r31 1 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.0900
+ $X2=0.5130 $Y2=0.0900
r32 10 21 0.314665 $w=2.27e-07 $l=4.5e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5130 $Y2=0.0900
.ends

.subckt PM_DFFLQNx3_ASAP7_75t_R%noxref_29 VSS 1
c1 1 VSS 0.00530465f
.ends

.subckt PM_DFFLQNx3_ASAP7_75t_R%SH VSS 11 12 13 14 78 81 86 89 17 25 27 15 6 18
+ 20 19 16 5 30 2 24 29 28 22 23 1 26 21
c1 1 VSS 0.00250926f
c2 2 VSS 0.0158733f
c3 5 VSS 0.00661763f
c4 6 VSS 0.00722138f
c5 11 VSS 0.0383819f
c6 12 VSS 0.0818527f
c7 13 VSS 0.0814081f
c8 14 VSS 0.081128f
c9 15 VSS 0.00490704f
c10 16 VSS 0.00512208f
c11 17 VSS 0.00843524f
c12 18 VSS 0.00193965f
c13 19 VSS 0.00224933f
c14 20 VSS 0.0025169f
c15 21 VSS 0.00125415f
c16 22 VSS 0.00137557f
c17 23 VSS 0.00250598f
c18 24 VSS 0.00429601f
c19 25 VSS 0.00657433f
c20 26 VSS 0.00318008f
c21 27 VSS 0.00102034f
c22 28 VSS 0.00123542f
c23 29 VSS 0.00117309f
c24 30 VSS 0.00358618f
r1 89 88 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r2 5 88 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6500 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r3 85 5 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6380 $Y=0.0405 $X2=0.6500 $Y2=0.0405
r4 15 85 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0405 $X2=0.6380 $Y2=0.0405
r5 86 15 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.0405 $X2=0.6335 $Y2=0.0405
r6 14 73 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=1.1070
+ $Y=0.1350 $X2=1.1070 $Y2=0.1360
r7 13 67 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=1.0530
+ $Y=0.1350 $X2=1.0530 $Y2=0.1360
r8 12 59 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.9990 $Y=0.1350 $X2=0.9990 $Y2=0.1360
r9 81 80 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r10 79 80 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7120 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r11 6 79 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7000 $Y=0.2295 $X2=0.7120 $Y2=0.2295
r12 16 6 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.2295 $X2=0.7000 $Y2=0.2295
r13 78 16 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.2295 $X2=0.6875 $Y2=0.2295
r14 5 57 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.0405
+ $X2=0.6480 $Y2=0.0360
r15 71 73 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.0945 $Y=0.1360 $X2=1.1070 $Y2=0.1360
r16 70 71 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.0800 $Y=0.1360 $X2=1.0945 $Y2=0.1360
r17 68 70 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.0655 $Y=0.1360 $X2=1.0800 $Y2=0.1360
r18 67 68 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.0530 $Y=0.1360 $X2=1.0655 $Y2=0.1360
r19 65 67 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.0405 $Y=0.1360 $X2=1.0530 $Y2=0.1360
r20 64 65 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.0260 $Y=0.1360 $X2=1.0405 $Y2=0.1360
r21 62 64 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.0115 $Y=0.1360 $X2=1.0260 $Y2=0.1360
r22 60 62 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=1.0085 $Y=0.1360 $X2=1.0115 $Y2=0.1360
r23 59 60 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.9990
+ $Y=0.1360 $X2=1.0085 $Y2=0.1360
r24 2 59 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.9895
+ $Y=0.1360 $X2=0.9990 $Y2=0.1360
r25 6 50 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7020 $Y=0.2295
+ $X2=0.7020 $Y2=0.2340
r26 57 58 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6480
+ $Y=0.0360 $X2=0.6615 $Y2=0.0360
r27 55 58 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0360 $X2=0.6615 $Y2=0.0360
r28 54 55 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6860
+ $Y=0.0360 $X2=0.6750 $Y2=0.0360
r29 17 26 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.7040
+ $Y=0.0360 $X2=0.7290 $Y2=0.0360
r30 17 54 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7040
+ $Y=0.0360 $X2=0.6860 $Y2=0.0360
r31 52 59 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.9990 $Y=0.1445
+ $X2=0.9990 $Y2=0.1360
r32 24 52 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.9990
+ $Y=0.1085 $X2=0.9990 $Y2=0.1445
r33 50 51 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.2340 $X2=0.7155 $Y2=0.2340
r34 25 51 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.2340 $X2=0.7155 $Y2=0.2340
r35 26 43 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.0360 $X2=0.7290 $Y2=0.0630
r36 47 52 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.9990 $Y=0.1530
+ $X2=0.9990 $Y2=0.1445
r37 46 47 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1530 $X2=0.9990 $Y2=0.1530
r38 45 46 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1530 $X2=0.9450 $Y2=0.1530
r39 30 45 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.8795
+ $Y=0.1530 $X2=0.8910 $Y2=0.1530
r40 44 45 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.8910 $Y=0.1485 $X2=0.8910
+ $Y2=0.1530
r41 23 44 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1305 $X2=0.8910 $Y2=0.1485
r42 19 39 6.50021 $w=1.33448e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1980 $X2=0.7290 $Y2=0.1690
r43 19 25 7.21452 $w=1.425e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1980 $X2=0.7290 $Y2=0.2340
r44 42 43 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.0900 $X2=0.7290 $Y2=0.0630
r45 41 42 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1090 $X2=0.7290 $Y2=0.0900
r46 18 27 4.67854 $w=1.44583e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1360 $X2=0.7290 $Y2=0.1600
r47 18 41 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1360 $X2=0.7290 $Y2=0.1090
r48 29 40 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1575 $X2=0.8910 $Y2=0.1665
r49 29 44 1.50855 $w=1.55e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1575 $X2=0.8910 $Y2=0.1485
r50 29 45 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.8910 $Y=0.1575 $X2=0.8910
+ $Y2=0.1530
r51 27 39 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1600 $X2=0.7290 $Y2=0.1690
r52 38 40 4.19024 $w=1.156e-08 $l=2.54018e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8660 $Y=0.1620 $X2=0.8910 $Y2=0.1665
r53 22 28 1.38478 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8480 $Y=0.1620 $X2=0.8370 $Y2=0.1620
r54 22 38 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8480
+ $Y=0.1620 $X2=0.8660 $Y2=0.1620
r55 37 39 4.4015 $w=1.35e-08 $l=2.78927e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7560 $Y=0.1620 $X2=0.7290 $Y2=0.1690
r56 36 37 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1620 $X2=0.7560 $Y2=0.1620
r57 20 28 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.1620 $X2=0.8370 $Y2=0.1620
r58 20 36 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.1620 $X2=0.7830 $Y2=0.1620
r59 28 35 4.88263 $w=1.47308e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8370 $Y=0.1620 $X2=0.8370 $Y2=0.1360
r60 21 35 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1180 $X2=0.8370 $Y2=0.1360
r61 34 35 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8370 $Y=0.1355
+ $X2=0.8370 $Y2=0.1360
r62 11 1 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.8370 $Y=0.1350 $X2=0.8370 $Y2=0.1245
r63 1 34 6.49795 $w=1.53e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08 $X=0.8370
+ $Y=0.1245 $X2=0.8370 $Y2=0.1355
.ends

.subckt PM_DFFLQNx3_ASAP7_75t_R%CLKB VSS 11 12 57 59 17 6 5 16 15 13 21 22 14
+ 19 18 2 1 20
c1 1 VSS 4.23044e-20
c2 2 VSS 0.000173057f
c3 5 VSS 0.00727948f
c4 6 VSS 0.00729137f
c5 11 VSS 0.00437566f
c6 12 VSS 0.0045835f
c7 13 VSS 0.00647745f
c8 14 VSS 0.00648564f
c9 15 VSS 0.0102281f
c10 16 VSS 0.00855722f
c11 17 VSS 0.00621822f
c12 18 VSS 0.000545754f
c13 19 VSS 0.00148618f
c14 20 VSS 0.00361003f
c15 21 VSS 0.00300575f
c16 22 VSS 0.0163679f
r1 14 6 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1600 $Y2=0.2160
r2 59 14 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r3 13 5 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1600 $Y2=0.0540
r4 57 13 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r5 6 53 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r6 5 50 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r7 53 54 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1845 $Y2=0.2340
r8 16 21 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.2340 $X2=0.2430 $Y2=0.2340
r9 16 54 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.1845 $Y2=0.2340
r10 50 51 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1845 $Y2=0.0360
r11 15 20 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.0360 $X2=0.2430 $Y2=0.0360
r12 15 51 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.1845 $Y2=0.0360
r13 2 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6750 $Y=0.1350
+ $X2=0.6750 $Y2=0.1440
r14 12 2 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6750
+ $Y=0.1350 $X2=0.6750 $Y2=0.1350
r15 21 44 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.2340 $X2=0.2430 $Y2=0.2125
r16 20 41 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0360 $X2=0.2430 $Y2=0.0575
r17 19 45 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1125 $X2=0.6750 $Y2=0.1440
r18 43 44 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1990 $X2=0.2430 $Y2=0.2125
r19 42 43 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1890 $X2=0.2430 $Y2=0.1990
r20 40 41 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0880 $X2=0.2430 $Y2=0.0575
r21 39 40 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1160 $X2=0.2430 $Y2=0.0880
r22 38 42 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1710 $X2=0.2430 $Y2=0.1890
r23 37 38 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1530 $X2=0.2430 $Y2=0.1710
r24 17 37 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1530
r25 17 39 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1160
r26 35 45 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.6750 $Y=0.1530
+ $X2=0.6750 $Y2=0.1440
r27 34 35 18.3054 $w=1.3e-08 $l=7.85e-08 $layer=M2 $thickness=3.6e-08 $X=0.5965
+ $Y=0.1530 $X2=0.6750 $Y2=0.1530
r28 33 34 29.3819 $w=1.3e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.4705
+ $Y=0.1530 $X2=0.5965 $Y2=0.1530
r29 32 33 15.2739 $w=1.3e-08 $l=6.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1530 $X2=0.4705 $Y2=0.1530
r30 31 32 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1530 $X2=0.4050 $Y2=0.1530
r31 30 31 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1530 $X2=0.3240 $Y2=0.1530
r32 30 37 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.2430 $Y=0.1530
+ $X2=0.2430 $Y2=0.1530
r33 22 30 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.2315
+ $Y=0.1530 $X2=0.2430 $Y2=0.1530
r34 28 32 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4050 $Y=0.1440
+ $X2=0.4050 $Y2=0.1530
r35 18 28 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1160 $X2=0.4050 $Y2=0.1440
r36 11 1 5.63117 $w=1.26721e-07 $l=2e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4050 $Y2=0.1330
r37 1 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1330
+ $X2=0.4050 $Y2=0.1440
.ends


*
.SUBCKT DFFLQNx3_ASAP7_75t_R VSS VDD CLK D QN
*
* VSS VSS
* VDD VDD
* CLK CLK
* D D
* QN QN
*
*

MM0 N_MM0_d N_MM0_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM27 N_MM27_d N_MM26_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM10_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM6 N_MM6_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM12 N_MM12_d N_MM12_g N_MM12_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM17 N_MM17_d N_MM13_g N_MM17_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM16 N_MM16_d N_MM19_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM14 N_MM14_d N_MM14_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM24 N_MM24_d N_MM24_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@3 N_MM24@3_d N_MM24@3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@2 N_MM24@2_d N_MM24@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM26 N_MM26_d N_MM26_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM13 N_MM13_d N_MM13_g N_MM13_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM18 N_MM18_d N_MM18_g N_MM18_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM19 N_MM19_d N_MM19_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM15 N_MM15_d N_MM14_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM25 N_MM25_d N_MM24_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@3 N_MM25@3_d N_MM24@3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@2 N_MM25@2_d N_MM24@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "DFFLQNx3_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "DFFLQNx3_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_DFFLQNx3_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_DFFLQNx3_ASAP7_75t_R%noxref_23
cc_1 N_noxref_23_1 N_MM3_g 0.0013737f
cc_2 N_noxref_23_1 N_CLKB_14 0.000769499f
cc_3 N_noxref_23_1 N_noxref_20_1 0.000469296f
cc_4 N_noxref_23_1 N_noxref_21_1 0.0076987f
cc_5 N_noxref_23_1 N_noxref_22_1 0.00123464f
x_PM_DFFLQNx3_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_DFFLQNx3_ASAP7_75t_R%noxref_22
cc_6 N_noxref_22_1 N_MM3_g 0.00136601f
cc_7 N_noxref_22_1 N_CLKB_13 0.0008021f
cc_8 N_noxref_22_1 N_noxref_20_1 0.00770196f
cc_9 N_noxref_22_1 N_noxref_21_1 0.000472628f
x_PM_DFFLQNx3_ASAP7_75t_R%PD4 VSS N_MM18_s N_MM19_d N_PD4_1
+ PM_DFFLQNx3_ASAP7_75t_R%PD4
cc_10 N_PD4_1 N_MM18_g 0.00773051f
cc_11 N_PD4_1 N_MM19_g 0.00776247f
x_PM_DFFLQNx3_ASAP7_75t_R%PD3 VSS N_MM9_s N_MM8_d N_PD3_1
+ PM_DFFLQNx3_ASAP7_75t_R%PD3
cc_12 N_PD3_1 N_MM9_g 0.00772309f
cc_13 N_PD3_1 N_MM11_g 0.00772966f
x_PM_DFFLQNx3_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_DFFLQNx3_ASAP7_75t_R%noxref_18
cc_14 N_noxref_18_1 N_MM0_g 0.00368932f
cc_15 N_noxref_18_1 N_CLKN_8 0.000543714f
cc_16 N_noxref_18_1 N_CLKN_9 4.21487e-20
cc_17 N_noxref_18_1 N_CLKN_31 5.87317e-20
cc_18 N_noxref_18_1 N_CLKN_23 0.000384559f
cc_19 N_noxref_18_1 N_CLKN_21 0.0276294f
x_PM_DFFLQNx3_ASAP7_75t_R%PU1 VSS N_MM3_d N_MM1_s N_PU1_1
+ PM_DFFLQNx3_ASAP7_75t_R%PU1
cc_20 N_PU1_1 N_MM1_g 0.0169384f
cc_21 N_PU1_1 N_MM3_g 0.0170113f
x_PM_DFFLQNx3_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_DFFLQNx3_ASAP7_75t_R%noxref_19
cc_22 N_noxref_19_1 N_MM0_g 0.00367453f
cc_23 N_noxref_19_1 N_CLKN_8 4.38676e-20
cc_24 N_noxref_19_1 N_CLKN_33 5.38656e-20
cc_25 N_noxref_19_1 N_CLKN_24 8.26328e-20
cc_26 N_noxref_19_1 N_CLKN_32 8.8491e-20
cc_27 N_noxref_19_1 N_CLKN_23 0.000271865f
cc_28 N_noxref_19_1 N_CLKN_9 0.00050327f
cc_29 N_noxref_19_1 N_CLKN_22 0.0277396f
cc_30 N_noxref_19_1 N_noxref_18_1 0.00204784f
x_PM_DFFLQNx3_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_DFFLQNx3_ASAP7_75t_R%noxref_21
cc_31 N_noxref_21_1 N_CLKN_1 0.000125863f
cc_32 N_noxref_21_1 N_MM26_g 0.00366742f
cc_33 N_noxref_21_1 N_CLKB_6 0.000435904f
cc_34 N_noxref_21_1 N_CLKB_14 0.0270926f
cc_35 N_noxref_21_1 N_noxref_20_1 0.00146986f
x_PM_DFFLQNx3_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_DFFLQNx3_ASAP7_75t_R%noxref_20
cc_36 N_noxref_20_1 N_CLKN_1 0.000129137f
cc_37 N_noxref_20_1 N_MM26_g 0.00352737f
cc_38 N_noxref_20_1 N_CLKB_5 0.000443316f
cc_39 N_noxref_20_1 N_CLKB_13 0.0271646f
x_PM_DFFLQNx3_ASAP7_75t_R%PD2 VSS N_MM10_s N_MM11_d N_PD2_5 N_PD2_1 N_PD2_4
+ PM_DFFLQNx3_ASAP7_75t_R%PD2
cc_40 N_PD2_5 N_CLKN_10 0.00146263f
cc_41 N_PD2_1 N_CLKN_3 0.00052085f
cc_42 N_PD2_1 N_MM9_g 0.00206401f
cc_43 N_PD2_4 N_MM9_g 0.00714445f
cc_44 N_PD2_5 N_MM9_g 0.0240626f
cc_45 N_PD2_4 N_MM10_g 0.0150104f
cc_46 N_PD2_5 N_MM11_g 0.0145937f
cc_47 N_PD2_1 N_MH_16 0.000461869f
cc_48 N_PD2_4 N_MH_3 0.000601242f
cc_49 N_PD2_1 N_MH_20 0.00323624f
x_PM_DFFLQNx3_ASAP7_75t_R%PD1 VSS N_MM5_d N_MM4_s N_PD1_5 N_PD1_4 N_PD1_1
+ PM_DFFLQNx3_ASAP7_75t_R%PD1
cc_50 N_PD1_5 N_CLKN_29 0.000206769f
cc_51 N_PD1_5 N_CLKN_2 0.00209484f
cc_52 N_PD1_5 N_MM1_g 0.073298f
cc_53 N_PD1_4 N_D_1 0.000671204f
cc_54 N_PD1_4 N_D_4 0.00076383f
cc_55 N_PD1_4 N_MM3_g 0.0361912f
cc_56 N_PD1_5 N_CLKB_18 0.000306124f
cc_57 N_PD1_5 N_CLKB_1 0.000757282f
cc_58 N_PD1_5 N_MM10_g 0.0346068f
cc_59 N_PD1_1 N_MH_4 0.00121055f
cc_60 N_PD1_1 N_MH_10 0.00348781f
x_PM_DFFLQNx3_ASAP7_75t_R%D VSS D N_MM3_g N_D_4 N_D_1 N_D_6 N_D_5
+ PM_DFFLQNx3_ASAP7_75t_R%D
cc_61 N_MM3_g N_CLKN_29 0.000914141f
cc_62 N_D_4 N_CLKN_36 0.000958413f
cc_63 N_D_1 N_CLKN_2 0.00239967f
cc_64 N_D_4 N_CLKN_29 0.00461049f
cc_65 N_MM3_g N_MM1_g 0.00524777f
x_PM_DFFLQNx3_ASAP7_75t_R%CLK VSS CLK N_MM0_g N_CLK_8 N_CLK_5 N_CLK_1 N_CLK_6
+ N_CLK_7 N_CLK_4 PM_DFFLQNx3_ASAP7_75t_R%CLK
x_PM_DFFLQNx3_ASAP7_75t_R%MH VSS N_MM7_g N_MM4_d N_MM9_d N_MM1_d N_MM10_d
+ N_MH_10 N_MH_20 N_MH_3 N_MH_16 N_MH_1 N_MH_17 N_MH_4 N_MH_12 N_MH_14 N_MH_18
+ N_MH_15 N_MH_19 PM_DFFLQNx3_ASAP7_75t_R%MH
cc_66 N_MH_10 N_CLKN_30 0.000373804f
cc_67 N_MH_10 N_MM1_g 0.000402462f
cc_68 N_MH_10 N_CLKN_29 0.000392264f
cc_69 N_MH_20 N_CLKN_30 0.000254848f
cc_70 N_MH_3 N_CLKN_2 0.000280463f
cc_71 N_MH_16 N_CLKN_30 0.00268685f
cc_72 N_MH_1 N_CLKN_10 0.00208808f
cc_73 N_MH_17 N_CLKN_10 0.000621088f
cc_74 N_MH_4 N_MM9_g 0.00063185f
cc_75 N_MH_16 N_CLKN_3 0.00076354f
cc_76 N_MH_12 N_CLKN_2 0.000880774f
cc_77 N_MH_3 N_CLKN_29 0.00133151f
cc_78 N_MH_14 N_CLKN_29 0.00140481f
cc_79 N_MH_14 N_CLKN_36 0.00151644f
cc_80 N_MH_3 N_MM1_g 0.00177588f
cc_81 N_MH_17 N_CLKN_30 0.00361758f
cc_82 N_MM7_g N_CLKN_10 0.00460022f
cc_83 N_MH_12 N_MM1_g 0.0337012f
cc_84 N_MM7_g N_MM12_g 0.0127509f
cc_85 N_MH_10 N_MM9_g 0.0363191f
cc_86 N_MH_10 N_MM13_g 0.00016165f
cc_87 N_MH_10 N_CLKB_18 0.000266086f
cc_88 N_MH_14 N_CLKB_18 0.000329917f
cc_89 N_MH_18 N_CLKB_18 0.000380679f
cc_90 N_MH_12 N_MM10_g 0.0164227f
cc_91 N_MH_3 N_CLKB_1 0.000736245f
cc_92 N_MH_4 N_MM10_g 0.00109537f
cc_93 N_MH_15 N_CLKB_18 0.00111834f
cc_94 N_MH_3 N_MM10_g 0.00117402f
cc_95 N_MH_17 N_CLKB_22 0.00124923f
cc_96 N_MH_16 N_CLKB_18 0.00135173f
cc_97 N_MH_12 N_CLKB_1 0.00182516f
cc_98 N_MH_16 N_CLKB_22 0.00225646f
cc_99 N_MH_19 N_CLKB_18 0.00273134f
cc_100 N_MH_10 N_MM10_g 0.0530825f
cc_101 N_MH_4 N_MS_1 0.000401778f
cc_102 N_MH_17 N_MS_18 0.000564021f
cc_103 N_MH_17 N_MS_1 0.000830126f
cc_104 N_MH_1 N_MS_14 0.000836332f
cc_105 N_MM7_g N_MS_3 0.000974805f
cc_106 N_MH_17 N_MS_17 0.00100383f
cc_107 N_MH_1 N_MM11_g 0.00106073f
cc_108 N_MM7_g N_MS_1 0.0011609f
cc_109 N_MH_15 N_MS_14 0.00123997f
cc_110 N_MM7_g N_MS_12 0.00639601f
cc_111 N_MM7_g N_MS_11 0.00640926f
cc_112 N_MH_17 N_MS_14 0.00719473f
cc_113 N_MM7_g N_MM11_g 0.0293056f
x_PM_DFFLQNx3_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_DFFLQNx3_ASAP7_75t_R%noxref_24
cc_114 N_noxref_24_1 N_SS_10 0.0170421f
cc_115 N_noxref_24_1 N_SH_1 0.00018406f
cc_116 N_noxref_24_1 N_MM14_g 0.0059476f
x_PM_DFFLQNx3_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_DFFLQNx3_ASAP7_75t_R%noxref_25
cc_117 N_noxref_25_1 N_SS_11 0.0168846f
cc_118 N_noxref_25_1 N_SH_1 0.000168104f
cc_119 N_noxref_25_1 N_MM14_g 0.00603655f
cc_120 N_noxref_25_1 N_noxref_24_1 0.00153921f
x_PM_DFFLQNx3_ASAP7_75t_R%SS VSS N_MM19_g N_MM14_d N_MM15_d N_SS_12 N_SS_10
+ N_SS_11 N_SS_4 N_SS_15 N_SS_3 N_SS_14 N_SS_1 N_SS_16 N_SS_13
+ PM_DFFLQNx3_ASAP7_75t_R%SS
cc_121 N_MM19_g N_CLKN_10 0.000218803f
cc_122 N_MM19_g N_CLKN_5 0.000537557f
cc_123 N_MM19_g N_MM18_g 0.0135466f
x_PM_DFFLQNx3_ASAP7_75t_R%PD5 VSS N_MM17_s N_MM16_d N_PD5_1 N_PD5_4 N_PD5_5
+ PM_DFFLQNx3_ASAP7_75t_R%PD5
cc_124 N_PD5_1 N_MM18_g 0.000859328f
cc_125 N_PD5_4 N_MM18_g 0.00695697f
cc_126 N_PD5_5 N_MM18_g 0.0239966f
cc_127 N_PD5_4 N_MM13_g 0.0152989f
cc_128 N_PD5_1 N_MM19_g 0.000917593f
cc_129 N_PD5_5 N_MM19_g 0.0155869f
cc_130 N_PD5_1 N_SH_15 0.000516331f
cc_131 N_PD5_1 N_SH_17 0.000458184f
cc_132 N_PD5_1 N_SH_18 0.000600155f
cc_133 N_PD5_4 N_SH_5 0.000661755f
cc_134 N_PD5_1 N_SH_26 0.00237749f
x_PM_DFFLQNx3_ASAP7_75t_R%noxref_28 VSS N_noxref_28_1
+ PM_DFFLQNx3_ASAP7_75t_R%noxref_28
cc_135 N_noxref_28_1 N_MM24@2_g 0.00147544f
cc_136 N_noxref_28_1 N_QN_14 0.037595f
x_PM_DFFLQNx3_ASAP7_75t_R%noxref_26 VSS N_noxref_26_1
+ PM_DFFLQNx3_ASAP7_75t_R%noxref_26
cc_137 N_noxref_26_1 N_SS_10 0.000650594f
cc_138 N_noxref_26_1 N_MM24_g 0.00172586f
cc_139 N_noxref_26_1 N_noxref_24_1 0.00775918f
cc_140 N_noxref_26_1 N_noxref_25_1 0.000476691f
x_PM_DFFLQNx3_ASAP7_75t_R%noxref_27 VSS N_noxref_27_1
+ PM_DFFLQNx3_ASAP7_75t_R%noxref_27
cc_141 N_noxref_27_1 N_SS_11 0.000640923f
cc_142 N_noxref_27_1 N_MM24_g 0.00173728f
cc_143 N_noxref_27_1 N_noxref_24_1 0.000478084f
cc_144 N_noxref_27_1 N_noxref_25_1 0.00775933f
cc_145 N_noxref_27_1 N_noxref_26_1 0.0012401f
x_PM_DFFLQNx3_ASAP7_75t_R%QN VSS QN N_MM24_d N_MM24@3_d N_MM24@2_d N_MM25_d
+ N_MM25@3_d N_MM25@2_d N_QN_13 N_QN_19 N_QN_18 N_QN_15 N_QN_3 N_QN_4 N_QN_1
+ N_QN_2 N_QN_16 N_QN_14 PM_DFFLQNx3_ASAP7_75t_R%QN
cc_146 N_QN_13 N_SH_24 0.00115571f
cc_147 N_QN_13 N_MM24@2_g 0.000884308f
cc_148 N_QN_13 N_SH_2 0.000468627f
cc_149 N_QN_13 N_SH_30 0.000715121f
cc_150 N_QN_19 N_SH_2 0.000819653f
cc_151 N_QN_18 N_MM24@2_g 0.000836474f
cc_152 N_QN_15 N_MM24@3_g 0.0308485f
cc_153 N_QN_3 N_MM24@2_g 0.000877682f
cc_154 N_QN_4 N_MM24@2_g 0.000941395f
cc_155 N_QN_1 N_SH_24 0.00155565f
cc_156 N_QN_1 N_MM24@3_g 0.00216426f
cc_157 N_QN_2 N_MM24@3_g 0.00218872f
cc_158 N_QN_16 N_MM24@2_g 0.0151636f
cc_159 N_QN_15 N_SH_2 0.00700132f
cc_160 N_QN_14 N_MM24@2_g 0.0524665f
cc_161 N_QN_13 N_MM24_g 0.0371148f
cc_162 N_QN_13 N_MM24@3_g 0.0683916f
x_PM_DFFLQNx3_ASAP7_75t_R%CLKN VSS N_MM26_g N_MM1_g N_MM9_g N_MM12_g N_MM18_g
+ N_MM0_d N_MM2_d N_CLKN_28 N_CLKN_35 N_CLKN_32 N_CLKN_9 N_CLKN_34 N_CLKN_8
+ N_CLKN_21 N_CLKN_22 N_CLKN_26 N_CLKN_25 N_CLKN_1 N_CLKN_27 N_CLKN_36
+ N_CLKN_23 N_CLKN_29 N_CLKN_2 N_CLKN_5 N_CLKN_30 N_CLKN_3 N_CLKN_10 N_CLKN_31
+ N_CLKN_33 N_CLKN_24 PM_DFFLQNx3_ASAP7_75t_R%CLKN
cc_163 N_CLKN_28 N_MM0_g 8.64818e-20
cc_164 N_CLKN_35 N_MM0_g 8.69563e-20
cc_165 N_CLKN_32 N_MM0_g 0.000192632f
cc_166 N_CLKN_9 N_MM0_g 0.00109915f
cc_167 N_CLKN_34 N_MM0_g 0.000233607f
cc_168 N_CLKN_8 N_MM0_g 0.00117509f
cc_169 N_CLKN_21 N_MM0_g 0.0112203f
cc_170 N_CLKN_22 N_MM0_g 0.0113257f
cc_171 N_CLKN_26 N_CLK_8 0.000734123f
cc_172 N_CLKN_25 N_CLK_5 0.000758513f
cc_173 N_CLKN_1 N_CLK_8 0.000777867f
cc_174 N_CLKN_27 N_CLK_1 0.000922771f
cc_175 N_CLKN_26 N_CLK_6 0.00131231f
cc_176 N_CLKN_27 N_CLK_7 0.00136568f
cc_177 N_CLKN_36 N_CLK_8 0.00169535f
cc_178 N_CLKN_23 N_CLK_4 0.00175957f
cc_179 N_CLKN_27 N_CLK_4 0.00214909f
cc_180 N_CLKN_34 N_CLK_8 0.00227131f
cc_181 N_CLKN_25 N_CLK_7 0.00227493f
cc_182 N_CLKN_1 N_CLK_1 0.00232584f
cc_183 N_CLKN_27 N_CLK_8 0.00241801f
cc_184 N_CLKN_32 N_CLK_8 0.00279116f
cc_185 N_MM26_g N_MM0_g 0.0351395f
x_PM_DFFLQNx3_ASAP7_75t_R%MS VSS N_MM11_g N_MM6_d N_MM12_d N_MM7_d N_MM13_d
+ N_MS_3 N_MS_11 N_MS_12 N_MS_13 N_MS_15 N_MS_1 N_MS_17 N_MS_4 N_MS_18 N_MS_14
+ N_MS_16 PM_DFFLQNx3_ASAP7_75t_R%MS
cc_186 N_MS_3 N_CLKN_30 0.000491949f
cc_187 N_MS_3 N_CLKN_10 0.000583097f
cc_188 N_MS_3 N_CLKN_3 0.000124014f
cc_189 N_MS_3 N_MM9_g 0.000162246f
cc_190 N_MS_3 N_CLKN_36 0.000188206f
cc_191 N_MS_11 N_MM12_g 0.00678254f
cc_192 N_MS_12 N_MM12_g 0.00780139f
cc_193 N_MS_13 N_MM12_g 0.00777423f
cc_194 N_MS_15 N_CLKN_10 0.000375043f
cc_195 N_MS_1 N_MM9_g 0.000568447f
cc_196 N_MS_17 N_CLKN_10 0.00155489f
cc_197 N_MS_4 N_MM12_g 0.00231983f
cc_198 N_MS_4 N_CLKN_10 0.00634581f
cc_199 N_MM11_g N_MM9_g 0.014383f
cc_200 N_MS_3 N_MM12_g 0.0257261f
cc_201 N_MS_13 N_MM10_g 0.000130191f
cc_202 N_MS_13 N_CLKB_19 0.00037352f
cc_203 N_MS_13 N_CLKB_22 0.000205471f
cc_204 N_MS_13 N_CLKB_2 0.000228055f
cc_205 N_MS_17 N_CLKB_19 0.00440571f
cc_206 N_MS_17 N_CLKB_2 0.00038569f
cc_207 N_MS_18 N_CLKB_19 0.000664924f
cc_208 N_MS_14 N_CLKB_22 0.00266996f
cc_209 N_MS_13 N_MM13_g 0.015394f
x_PM_DFFLQNx3_ASAP7_75t_R%noxref_29 VSS N_noxref_29_1
+ PM_DFFLQNx3_ASAP7_75t_R%noxref_29
cc_210 N_noxref_29_1 N_MM24@2_g 0.00147935f
cc_211 N_noxref_29_1 N_QN_16 0.0378692f
cc_212 N_noxref_29_1 N_noxref_28_1 0.00176738f
x_PM_DFFLQNx3_ASAP7_75t_R%SH VSS N_MM14_g N_MM24_g N_MM24@3_g N_MM24@2_g
+ N_MM13_s N_MM18_d N_MM12_s N_MM17_d N_SH_17 N_SH_25 N_SH_27 N_SH_15 N_SH_6
+ N_SH_18 N_SH_20 N_SH_19 N_SH_16 N_SH_5 N_SH_30 N_SH_2 N_SH_24 N_SH_29 N_SH_28
+ N_SH_22 N_SH_23 N_SH_1 N_SH_26 N_SH_21 PM_DFFLQNx3_ASAP7_75t_R%SH
cc_213 N_SH_17 N_CLKN_36 0.000109007f
cc_214 N_SH_25 N_CLKN_10 0.000173184f
cc_215 N_SH_27 N_CLKN_10 0.000204456f
cc_216 N_SH_15 N_MM12_g 0.00677846f
cc_217 N_SH_6 N_CLKN_10 0.000267105f
cc_218 N_SH_18 N_CLKN_10 0.000419691f
cc_219 N_SH_20 N_CLKN_5 0.000428302f
cc_220 N_SH_19 N_CLKN_10 0.000620804f
cc_221 N_SH_16 N_CLKN_5 0.000929177f
cc_222 N_SH_6 N_MM18_g 0.0010039f
cc_223 N_SH_16 N_CLKN_10 0.00226816f
cc_224 N_SH_5 N_MM12_g 0.00951821f
cc_225 N_SH_16 N_MM18_g 0.0162828f
cc_226 N_SH_30 N_CLKB_22 0.000137311f
cc_227 N_SH_6 N_MM13_g 0.000141727f
cc_228 N_SH_20 N_CLKB_19 0.000214028f
cc_229 N_SH_16 N_MM13_g 0.00675261f
cc_230 N_SH_15 N_MM13_g 0.00679213f
cc_231 N_SH_25 N_CLKB_19 0.0003116f
cc_232 N_SH_27 N_CLKB_19 0.00094534f
cc_233 N_SH_18 N_CLKB_2 0.000463902f
cc_234 N_SH_5 N_CLKB_2 0.000532303f
cc_235 N_SH_19 N_CLKB_19 0.000538342f
cc_236 N_SH_17 N_CLKB_19 0.000565326f
cc_237 N_SH_17 N_CLKB_22 0.00105009f
cc_238 N_SH_18 N_CLKB_19 0.00407762f
cc_239 N_SH_5 N_MM13_g 0.0184274f
cc_240 N_SH_19 N_MS_3 0.000109634f
cc_241 N_SH_18 N_MS_3 0.000116089f
cc_242 N_SH_25 N_MS_3 0.000158325f
cc_243 N_SH_16 N_MS_3 0.000437606f
cc_244 N_SH_15 N_MS_3 0.000465255f
cc_245 N_SH_6 N_MS_4 0.000686016f
cc_246 N_SH_25 N_MS_4 0.00029747f
cc_247 N_SH_25 N_MS_17 0.000539992f
cc_248 N_SH_17 N_MS_16 0.000589665f
cc_249 N_SH_16 N_MS_4 0.000599966f
cc_250 N_SH_17 N_MS_18 0.00163972f
cc_251 N_SH_5 N_MS_3 0.00362309f
cc_252 N_SH_17 N_MM19_g 0.000115713f
cc_253 N_SH_19 N_MM19_g 0.000128107f
cc_254 N_SH_2 N_MM19_g 0.000169893f
cc_255 N_SH_24 N_MM19_g 0.000175165f
cc_256 N_SH_29 N_MM19_g 0.000183487f
cc_257 N_SH_28 N_SS_12 0.000219151f
cc_258 N_MM14_g N_SS_10 0.00686385f
cc_259 N_MM14_g N_SS_11 0.00682884f
cc_260 N_SH_22 N_SS_4 0.000249496f
cc_261 N_SH_2 N_SS_15 0.00027392f
cc_262 N_SH_24 N_SS_15 0.00722616f
cc_263 N_MM14_g N_SS_3 0.000405f
cc_264 N_SH_23 N_SS_15 0.00188115f
cc_265 N_MM14_g N_SS_4 0.000527123f
cc_266 N_SH_22 N_SS_14 0.000651366f
cc_267 N_SH_1 N_SS_1 0.00070153f
cc_268 N_SH_26 N_SS_16 0.000793581f
cc_269 N_SH_18 N_SS_1 0.000844674f
cc_270 N_SH_29 N_SS_15 0.000900665f
cc_271 N_SH_21 N_SS_12 0.000937997f
cc_272 N_MM14_g N_SS_1 0.00110551f
cc_273 N_SH_23 N_SS_13 0.00110841f
cc_274 N_SH_1 N_MM19_g 0.00113664f
cc_275 N_SH_29 N_SS_14 0.00128222f
cc_276 N_SH_20 N_SS_12 0.00157249f
cc_277 N_SH_30 N_SS_15 0.00189009f
cc_278 N_SH_18 N_SS_12 0.00471933f
cc_279 N_MM14_g N_MM19_g 0.0293845f
x_PM_DFFLQNx3_ASAP7_75t_R%CLKB VSS N_MM10_g N_MM13_g N_MM27_d N_MM26_d
+ N_CLKB_17 N_CLKB_6 N_CLKB_5 N_CLKB_16 N_CLKB_15 N_CLKB_13 N_CLKB_21 N_CLKB_22
+ N_CLKB_14 N_CLKB_19 N_CLKB_18 N_CLKB_2 N_CLKB_1 N_CLKB_20
+ PM_DFFLQNx3_ASAP7_75t_R%CLKB
cc_280 N_CLKB_17 N_CLK_5 9.42652e-20
cc_281 N_CLKB_6 N_CLK_5 0.000321239f
cc_282 N_CLKB_5 N_CLK_5 0.000406233f
cc_283 N_CLKB_16 N_CLK_5 0.000213606f
cc_284 N_CLKB_16 N_CLK_6 0.000974336f
cc_285 N_CLKB_15 N_CLK_5 0.00222408f
cc_286 N_CLKB_13 N_CLKN_26 3.22363e-20
cc_287 N_CLKB_13 N_CLKN_23 6.63422e-20
cc_288 N_MM13_g N_CLKN_5 0.000222584f
cc_289 N_CLKB_21 N_CLKN_34 0.000231065f
cc_290 N_CLKB_6 N_CLKN_34 0.000271072f
cc_291 N_CLKB_22 N_CLKN_30 0.000665549f
cc_292 N_CLKB_6 N_CLKN_1 0.000308943f
cc_293 N_CLKB_14 N_MM26_g 0.0112471f
cc_294 N_CLKB_16 N_CLKN_34 0.00508495f
cc_295 N_CLKB_22 N_CLKN_29 0.000355479f
cc_296 N_CLKB_15 N_CLKN_35 0.000446f
cc_297 N_MM10_g N_CLKN_3 0.000540881f
cc_298 N_CLKB_19 N_CLKN_10 0.000573168f
cc_299 N_CLKB_18 N_CLKN_36 0.000611247f
cc_300 N_CLKB_14 N_CLKN_1 0.000622622f
cc_301 N_CLKB_6 N_CLKN_27 0.000664076f
cc_302 N_CLKB_2 N_CLKN_10 0.00285577f
cc_303 N_CLKB_17 N_CLKN_36 0.000735061f
cc_304 N_CLKB_5 N_MM26_g 0.000758246f
cc_305 N_CLKB_1 N_CLKN_2 0.00227225f
cc_306 N_CLKB_17 N_CLKN_28 0.000987161f
cc_307 N_CLKB_6 N_MM26_g 0.00107449f
cc_308 N_MM10_g N_MM1_g 0.0016279f
cc_309 N_CLKB_18 N_CLKN_29 0.00310318f
cc_310 N_CLKB_17 N_CLKN_35 0.00376576f
cc_311 N_MM13_g N_CLKN_10 0.00430634f
cc_312 N_MM13_g N_MM12_g 0.00567058f
cc_313 N_MM10_g N_MM9_g 0.00910719f
cc_314 N_MM13_g N_MM18_g 0.0184478f
cc_315 N_CLKB_22 N_CLKN_36 0.0282491f
cc_316 N_CLKB_13 N_MM26_g 0.038841f
cc_317 N_CLKB_18 N_D_4 0.000146015f
cc_318 N_CLKB_21 N_D_6 0.000777105f
cc_319 N_CLKB_20 N_D_5 0.00096655f
cc_320 N_CLKB_22 N_D_4 0.0010836f
cc_321 N_CLKB_17 N_D_4 0.00840269f
*END of DFFLQNx3_ASAP7_75t_R.pxi
.ENDS
** Design:	DFFLQx4_ASAP7_75t_R
* Created:	"Fri Aug 17 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "DFFLQx4_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "DFFLQx4_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_DFFLQx4_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.041829f
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.0418025f
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%noxref_29 VSS 1
c1 1 VSS 0.0422386f
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%noxref_30 VSS 1
c1 1 VSS 0.0422876f
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%Q VSS 35 26 27 41 42 50 51 54 55 14 18 16 15 13
+ 21 20 2 3 4 1
c1 1 VSS 0.00896245f
c2 2 VSS 0.00879007f
c3 3 VSS 0.00949353f
c4 4 VSS 0.0100404f
c5 13 VSS 0.00449484f
c6 14 VSS 0.00445184f
c7 15 VSS 0.00444822f
c8 16 VSS 0.00439491f
c9 17 VSS 0.0166987f
c10 18 VSS 0.0170306f
c11 19 VSS 0.00775942f
c12 20 VSS 0.00288773f
c13 21 VSS 0.00342659f
c14 22 VSS 0.00326813f
c15 23 VSS 0.00325127f
r1 55 53 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.1510 $Y=0.2025 $X2=1.1485 $Y2=0.2025
r2 2 53 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.1340 $Y=0.2025 $X2=1.1485 $Y2=0.2025
r3 15 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.1195 $Y=0.2025 $X2=1.1340 $Y2=0.2025
r4 54 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.1170 $Y=0.2025 $X2=1.1195 $Y2=0.2025
r5 2 47 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.1340 $Y=0.2025
+ $X2=1.1340 $Y2=0.2160
r6 51 49 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.2590 $Y=0.2025 $X2=1.2565 $Y2=0.2025
r7 4 49 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.2420 $Y=0.2025 $X2=1.2565 $Y2=0.2025
r8 16 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.2275 $Y=0.2025 $X2=1.2420 $Y2=0.2025
r9 50 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.2250 $Y=0.2025 $X2=1.2275 $Y2=0.2025
r10 21 45 4.64944 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.1340
+ $Y=0.2340 $X2=1.1590 $Y2=0.2340
r11 21 47 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.1340
+ $Y=0.2340 $X2=1.1340 $Y2=0.2160
r12 4 43 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.2420 $Y=0.2025
+ $X2=1.2420 $Y2=0.2340
r13 43 44 9.32759 $w=1.3e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=1.2420
+ $Y=0.2340 $X2=1.2820 $Y2=0.2340
r14 18 43 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.2040
+ $Y=0.2340 $X2=1.2420 $Y2=0.2340
r15 18 45 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.2040
+ $Y=0.2340 $X2=1.1590 $Y2=0.2340
r16 23 38 2.48126 $w=1.71429e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3230 $Y=0.2340 $X2=1.3230 $Y2=0.2130
r17 23 44 7.66726 $w=1.56829e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3230 $Y=0.2340 $X2=1.2820 $Y2=0.2340
r18 42 40 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.2590 $Y=0.0675 $X2=1.2565 $Y2=0.0675
r19 3 40 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.2420 $Y=0.0675 $X2=1.2565 $Y2=0.0675
r20 14 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.2275 $Y=0.0675 $X2=1.2420 $Y2=0.0675
r21 41 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.2250 $Y=0.0675 $X2=1.2275 $Y2=0.0675
r22 37 38 6.8096 $w=1.5e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.1730 $X2=1.3230 $Y2=0.2130
r23 36 37 5.66048 $w=1.5e-08 $l=3.33e-08 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.1397 $X2=1.3230 $Y2=0.1730
r24 35 36 0.97888 $w=1.5e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.1340 $X2=1.3230 $Y2=0.1397
r25 35 34 0.6384 $w=1.5e-08 $l=3.8e-09 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.1340 $X2=1.3230 $Y2=0.1302
r26 33 34 5.49024 $w=1.5e-08 $l=3.22e-08 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.0980 $X2=1.3230 $Y2=0.1302
r27 19 22 2.48126 $w=1.71429e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3230 $Y=0.0570 $X2=1.3230 $Y2=0.0360
r28 19 33 6.97984 $w=1.5e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.0570 $X2=1.3230 $Y2=0.0980
r29 3 31 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.2420 $Y=0.0675
+ $X2=1.2420 $Y2=0.0360
r30 22 32 7.66726 $w=1.56829e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3230 $Y=0.0360 $X2=1.2820 $Y2=0.0360
r31 31 32 9.32759 $w=1.3e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=1.2420
+ $Y=0.0360 $X2=1.2820 $Y2=0.0360
r32 30 31 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.2040
+ $Y=0.0360 $X2=1.2420 $Y2=0.0360
r33 17 29 4.64944 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.1590
+ $Y=0.0360 $X2=1.1340 $Y2=0.0360
r34 17 30 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.1590
+ $Y=0.0360 $X2=1.2040 $Y2=0.0360
r35 20 29 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.1340
+ $Y=0.0540 $X2=1.1340 $Y2=0.0360
r36 1 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.1340 $Y=0.0675
+ $X2=1.1340 $Y2=0.0540
r37 27 25 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.1510 $Y=0.0675 $X2=1.1485 $Y2=0.0675
r38 1 25 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.1340 $Y=0.0675 $X2=1.1485 $Y2=0.0675
r39 13 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.1195 $Y=0.0675 $X2=1.1340 $Y2=0.0675
r40 26 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.1170 $Y=0.0675 $X2=1.1195 $Y2=0.0675
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%noxref_28 VSS 1
c1 1 VSS 0.0415404f
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%noxref_26 VSS 1
c1 1 VSS 0.00423821f
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%QN VSS 9 10 11 12 62 63 66 67 13 16 4 17 18 14 3
+ 1 22 20 19
c1 1 VSS 0.0190282f
c2 3 VSS 0.013207f
c3 4 VSS 0.01375f
c4 9 VSS 0.0817182f
c5 10 VSS 0.0814426f
c6 11 VSS 0.0816427f
c7 12 VSS 0.0820944f
c8 13 VSS 0.00823584f
c9 14 VSS 0.00822929f
c10 15 VSS 0.00924858f
c11 16 VSS 0.00859447f
c12 17 VSS 0.00393659f
c13 18 VSS 0.00383258f
c14 19 VSS 0.00289309f
c15 20 VSS 0.00432824f
c16 21 VSS 0.00143057f
c17 22 VSS 0.00355558f
r1 67 65 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0430 $Y=0.2025 $X2=1.0405 $Y2=0.2025
r2 4 65 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0260 $Y=0.2025 $X2=1.0405 $Y2=0.2025
r3 14 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0115 $Y=0.2025 $X2=1.0260 $Y2=0.2025
r4 66 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0090 $Y=0.2025 $X2=1.0115 $Y2=0.2025
r5 63 61 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.0430 $Y=0.0675 $X2=1.0405 $Y2=0.0675
r6 3 61 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.0260 $Y=0.0675 $X2=1.0405 $Y2=0.0675
r7 13 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.0115 $Y=0.0675 $X2=1.0260 $Y2=0.0675
r8 62 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.0090 $Y=0.0675 $X2=1.0115 $Y2=0.0675
r9 4 58 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0260 $Y=0.2025
+ $X2=1.0260 $Y2=0.2340
r10 3 56 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0260 $Y=0.0675
+ $X2=1.0260 $Y2=0.0360
r11 58 59 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.2340 $X2=1.0575 $Y2=0.2340
r12 16 58 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.0145
+ $Y=0.2340 $X2=1.0260 $Y2=0.2340
r13 56 57 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.0360 $X2=1.0575 $Y2=0.0360
r14 15 56 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.0145
+ $Y=0.0360 $X2=1.0260 $Y2=0.0360
r15 22 55 3.24787 $w=1.72e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.0890
+ $Y=0.2340 $X2=1.0890 $Y2=0.2130
r16 22 59 5.69637 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0890 $Y=0.2340 $X2=1.0575 $Y2=0.2340
r17 20 53 3.24787 $w=1.72e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.0890
+ $Y=0.0360 $X2=1.0890 $Y2=0.0570
r18 20 57 5.69637 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0890 $Y=0.0360 $X2=1.0575 $Y2=0.0360
r19 54 55 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=1.0890
+ $Y=0.1840 $X2=1.0890 $Y2=0.2130
r20 18 21 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=1.0890
+ $Y=0.1560 $X2=1.0890 $Y2=0.1360
r21 18 54 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.0890
+ $Y=0.1560 $X2=1.0890 $Y2=0.1840
r22 52 53 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=1.0890
+ $Y=0.0955 $X2=1.0890 $Y2=0.0570
r23 17 21 1.50137 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0890 $Y=0.1245 $X2=1.0890 $Y2=0.1360
r24 17 52 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=1.0890
+ $Y=0.1245 $X2=1.0890 $Y2=0.0955
r25 21 49 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.0890
+ $Y=0.1360 $X2=1.1115 $Y2=0.1360
r26 12 43 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=1.2690
+ $Y=0.1350 $X2=1.2690 $Y2=0.1360
r27 11 37 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=1.2150
+ $Y=0.1350 $X2=1.2150 $Y2=0.1360
r28 48 49 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.1340
+ $Y=0.1360 $X2=1.1115 $Y2=0.1360
r29 19 46 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.1475
+ $Y=0.1360 $X2=1.1610 $Y2=0.1360
r30 19 48 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.1475
+ $Y=0.1360 $X2=1.1340 $Y2=0.1360
r31 10 30 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=1.1610 $Y=0.1350 $X2=1.1610 $Y2=0.1360
r32 41 43 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.2565 $Y=0.1360 $X2=1.2690 $Y2=0.1360
r33 40 41 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.2420 $Y=0.1360 $X2=1.2565 $Y2=0.1360
r34 38 40 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.2275 $Y=0.1360 $X2=1.2420 $Y2=0.1360
r35 37 38 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.2150 $Y=0.1360 $X2=1.2275 $Y2=0.1360
r36 35 37 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.2025 $Y=0.1360 $X2=1.2150 $Y2=0.1360
r37 34 35 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.1880 $Y=0.1360 $X2=1.2025 $Y2=0.1360
r38 32 34 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.1735 $Y=0.1360 $X2=1.1880 $Y2=0.1360
r39 31 32 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=1.1705 $Y=0.1360 $X2=1.1735 $Y2=0.1360
r40 30 31 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=1.1610
+ $Y=0.1360 $X2=1.1705 $Y2=0.1360
r41 30 46 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.1610 $Y=0.1360
+ $X2=1.1610 $Y2=0.1360
r42 29 30 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=1.1515
+ $Y=0.1360 $X2=1.1610 $Y2=0.1360
r43 27 29 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=1.1485 $Y=0.1360 $X2=1.1515 $Y2=0.1360
r44 26 27 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.1340 $Y=0.1360 $X2=1.1485 $Y2=0.1360
r45 25 26 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.1195 $Y=0.1360 $X2=1.1340 $Y2=0.1360
r46 9 1 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=1.1070
+ $Y=0.1350 $X2=1.1070 $Y2=0.1360
r47 1 24 2.90696 $w=2.1681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.1070 $Y=0.1360 $X2=1.0965 $Y2=0.1360
r48 1 25 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.1070 $Y=0.1360 $X2=1.1195 $Y2=0.1360
r49 9 24 0.610027 $w=2.16919e-07 $l=1.05475e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=1.1070 $Y=0.1350 $X2=1.0965 $Y2=0.1360
r50 9 25 1.79147 $w=1.8466e-07 $l=1.25399e-08 $layer=LIG $thickness=5.44e-08
+ $X=1.1070 $Y=0.1350 $X2=1.1195 $Y2=0.1360
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%noxref_27 VSS 1
c1 1 VSS 0.0415022f
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.00421443f
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%D VSS 9 3 1 4 6 5
c1 1 VSS 0.00689107f
c2 3 VSS 0.0834372f
c3 4 VSS 0.00587845f
c4 5 VSS 0.00710926f
c5 6 VSS 0.00759484f
r1 6 13 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.2340 $X2=0.2970 $Y2=0.2140
r2 5 8 5.17411 $w=1.46514e-08 $l=2.72e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0360 $X2=0.2970 $Y2=0.0632
r3 12 13 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1735 $X2=0.2970 $Y2=0.2140
r4 11 12 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1735
r5 9 10 2.85657 $w=1.3e-08 $l=1.22e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0820 $X2=0.2970 $Y2=0.0942
r6 9 8 4.37231 $w=1.3e-08 $l=1.88e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0820 $X2=0.2970 $Y2=0.0632
r7 4 10 5.07188 $w=1.3e-08 $l=2.18e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1160 $X2=0.2970 $Y2=0.0942
r8 4 11 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1160 $X2=0.2970 $Y2=0.1350
r9 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r10 1 11 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%CLK VSS 11 3 8 5 1 6 7 4
c1 1 VSS 0.00249851f
c2 3 VSS 0.0597519f
c3 4 VSS 0.000981185f
c4 5 VSS 0.00400902f
c5 6 VSS 0.00368869f
c6 7 VSS 0.00232012f
c7 8 VSS 0.00194789f
r1 6 17 3.22357 $w=2.26279e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.2125 $X2=0.1080 $Y2=0.1820
r2 5 15 3.22357 $w=2.26279e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0575 $X2=0.1080 $Y2=0.0880
r3 16 17 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.1820 $X2=0.1080 $Y2=0.1820
r4 8 13 2.6406 $w=2.38947e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1820 $X2=0.0810 $Y2=0.1540
r5 8 16 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1820 $X2=0.0945 $Y2=0.1820
r6 14 15 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.0880 $X2=0.1080 $Y2=0.0880
r7 7 10 1.76614 $w=2.65738e-08 $l=2.42e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0880 $X2=0.0810 $Y2=0.1122
r8 7 14 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0880 $X2=0.0945 $Y2=0.0880
r9 11 12 0.874462 $w=1.3e-08 $l=3.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1227
r10 11 10 1.57403 $w=1.3e-08 $l=6.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1122
r11 4 12 2.85657 $w=1.3e-08 $l=1.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1227
r12 4 13 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1540
r13 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r14 1 4 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%PD3 VSS 2 4 1
c1 1 VSS 0.000973923f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0405 $X2=0.4905 $Y2=0.0405
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0405 $X2=0.4735 $Y2=0.0405
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4735 $Y=0.0405 $X2=0.4905 $Y2=0.0405
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%PD2 VSS 7 12 4 1 5
c1 1 VSS 0.00724145f
c2 4 VSS 0.00187201f
c3 5 VSS 0.00234338f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4880 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r3 9 5 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.4605
+ $Y=0.2295 $X2=0.4860 $Y2=0.2295
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.4455
+ $Y=0.2295 $X2=0.4605 $Y2=0.2295
r5 1 8 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4320
+ $Y=0.2295 $X2=0.4455 $Y2=0.2295
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2295 $X2=0.4300 $Y2=0.2295
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2295 $X2=0.4175 $Y2=0.2295
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%PU1 VSS 2 4 1
c1 1 VSS 0.000978334f
r1 4 3 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3365 $Y2=0.2025
r2 2 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3195 $Y2=0.2025
r3 1 3 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3195 $Y=0.2025 $X2=0.3365 $Y2=0.2025
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%PD4 VSS 2 4 1
c1 1 VSS 0.000946814f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.2295 $X2=0.7605 $Y2=0.2295
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.2295 $X2=0.7435 $Y2=0.2295
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7435 $Y=0.2295 $X2=0.7605 $Y2=0.2295
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%MS VSS 10 39 42 47 49 3 15 13 12 1 17 11 4 18 14
+ 16
c1 1 VSS 0.00220354f
c2 3 VSS 0.00515006f
c3 4 VSS 0.00958327f
c4 10 VSS 0.0375403f
c5 11 VSS 0.00286534f
c6 12 VSS 0.00270673f
c7 13 VSS 0.00224998f
c8 14 VSS 0.00193957f
c9 15 VSS 0.00423155f
c10 16 VSS 0.00291708f
c11 17 VSS 0.00105151f
c12 18 VSS 0.000406705f
c13 19 VSS 0.00265754f
r1 49 48 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.2295 $X2=0.6625 $Y2=0.2295
r2 13 48 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6500 $Y=0.2295 $X2=0.6625 $Y2=0.2295
r3 12 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2295 $X2=0.5920 $Y2=0.2295
r4 47 12 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.2295 $X2=0.5795 $Y2=0.2295
r5 44 13 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6210 $Y=0.2295 $X2=0.6480 $Y2=0.2295
r6 4 44 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08 $X=0.5940
+ $Y=0.2295 $X2=0.6210 $Y2=0.2295
r7 4 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2295
+ $X2=0.5965 $Y2=0.2340
r8 15 19 4.06404 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5965 $Y=0.2340 $X2=0.6210 $Y2=0.2340
r9 42 41 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.0405 $X2=0.6085 $Y2=0.0405
r10 40 41 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6040 $Y=0.0405 $X2=0.6085 $Y2=0.0405
r11 3 40 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5920 $Y=0.0405 $X2=0.6040 $Y2=0.0405
r12 11 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.0405 $X2=0.5920 $Y2=0.0405
r13 39 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0405 $X2=0.5795 $Y2=0.0405
r14 19 35 3.01468 $w=1.741e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.2340 $X2=0.6210 $Y2=0.2140
r15 3 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0405
+ $X2=0.5940 $Y2=0.0540
r16 34 35 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1850 $X2=0.6210 $Y2=0.2140
r17 33 34 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1660 $X2=0.6210 $Y2=0.1850
r18 32 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1525 $X2=0.6210 $Y2=0.1660
r19 31 32 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1310 $X2=0.6210 $Y2=0.1525
r20 17 28 3.60008 $w=1.51951e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.1105 $X2=0.6210 $Y2=0.0900
r21 17 31 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1105 $X2=0.6210 $Y2=0.1310
r22 16 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0540 $X2=0.5940 $Y2=0.0720
r23 27 28 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6075 $Y=0.0900 $X2=0.6210 $Y2=0.0900
r24 18 26 1.38478 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5940 $Y=0.0900 $X2=0.5830 $Y2=0.0900
r25 18 27 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5940 $Y=0.0900 $X2=0.6075 $Y2=0.0900
r26 18 29 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0900 $X2=0.5940 $Y2=0.0720
r27 25 26 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5515
+ $Y=0.0900 $X2=0.5830 $Y2=0.0900
r28 24 25 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0900 $X2=0.5515 $Y2=0.0900
r29 14 24 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5000
+ $Y=0.0900 $X2=0.5130 $Y2=0.0900
r30 1 21 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.5130
+ $Y=0.0900 $X2=0.5130 $Y2=0.0900
r31 1 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.0900
+ $X2=0.5130 $Y2=0.0900
r32 10 21 0.314665 $w=2.27e-07 $l=4.5e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5130 $Y2=0.0900
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.00426358f
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.00474072f
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.00432266f
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%PD1 VSS 7 10 4 5 1
c1 1 VSS 0.00937213f
c2 4 VSS 0.00316343f
c3 5 VSS 0.00185665f
r1 10 9 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r2 8 9 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r3 5 8 0.123457 $w=8.1e-08 $l=1e-08 $layer=N_src_drn $thickness=1e-09 $X=0.3780
+ $Y=0.0675 $X2=0.3880 $Y2=0.0675
r4 4 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3220 $Y2=0.0675
r5 7 4 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r6 1 5 1e-05
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.00476662f
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%CLKB VSS 11 12 57 59 17 6 5 16 15 13 21 22 14 19
+ 18 2 1 20
c1 1 VSS 3.14663e-20
c2 2 VSS 0.00016845f
c3 5 VSS 0.0073337f
c4 6 VSS 0.00735435f
c5 11 VSS 0.00437749f
c6 12 VSS 0.00458025f
c7 13 VSS 0.00632813f
c8 14 VSS 0.0063526f
c9 15 VSS 0.00851004f
c10 16 VSS 0.00870945f
c11 17 VSS 0.00618853f
c12 18 VSS 0.000537921f
c13 19 VSS 0.00143342f
c14 20 VSS 0.00355513f
c15 21 VSS 0.00287596f
c16 22 VSS 0.0154922f
r1 14 6 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1600 $Y2=0.2160
r2 59 14 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r3 13 5 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1600 $Y2=0.0540
r4 57 13 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r5 6 53 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r6 5 50 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r7 53 54 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1845 $Y2=0.2340
r8 16 21 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.2340 $X2=0.2430 $Y2=0.2340
r9 16 54 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.1845 $Y2=0.2340
r10 50 51 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1845 $Y2=0.0360
r11 15 20 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.0360 $X2=0.2430 $Y2=0.0360
r12 15 51 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.1845 $Y2=0.0360
r13 2 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6750 $Y=0.1350
+ $X2=0.6750 $Y2=0.1440
r14 12 2 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6750
+ $Y=0.1350 $X2=0.6750 $Y2=0.1350
r15 21 44 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.2340 $X2=0.2430 $Y2=0.2125
r16 20 41 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0360 $X2=0.2430 $Y2=0.0575
r17 19 45 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1125 $X2=0.6750 $Y2=0.1440
r18 43 44 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1990 $X2=0.2430 $Y2=0.2125
r19 42 43 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1890 $X2=0.2430 $Y2=0.1990
r20 40 41 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0880 $X2=0.2430 $Y2=0.0575
r21 39 40 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1160 $X2=0.2430 $Y2=0.0880
r22 38 42 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1710 $X2=0.2430 $Y2=0.1890
r23 37 38 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1530 $X2=0.2430 $Y2=0.1710
r24 17 37 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1530
r25 17 39 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1160
r26 35 45 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.6750 $Y=0.1530
+ $X2=0.6750 $Y2=0.1440
r27 34 35 18.3054 $w=1.3e-08 $l=7.85e-08 $layer=M2 $thickness=3.6e-08 $X=0.5965
+ $Y=0.1530 $X2=0.6750 $Y2=0.1530
r28 33 34 29.3819 $w=1.3e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.4705
+ $Y=0.1530 $X2=0.5965 $Y2=0.1530
r29 32 33 15.2739 $w=1.3e-08 $l=6.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1530 $X2=0.4705 $Y2=0.1530
r30 31 32 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1530 $X2=0.4050 $Y2=0.1530
r31 30 31 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1530 $X2=0.3240 $Y2=0.1530
r32 30 37 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.2430 $Y=0.1530
+ $X2=0.2430 $Y2=0.1530
r33 22 30 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.2315
+ $Y=0.1530 $X2=0.2430 $Y2=0.1530
r34 28 32 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4050 $Y=0.1440
+ $X2=0.4050 $Y2=0.1530
r35 18 28 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1160 $X2=0.4050 $Y2=0.1440
r36 11 1 5.63117 $w=1.26721e-07 $l=2e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4050 $Y2=0.1330
r37 1 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1330
+ $X2=0.4050 $Y2=0.1440
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%PD5 VSS 7 12 1 5 4
c1 1 VSS 0.0074908f
c2 4 VSS 0.00188428f
c3 5 VSS 0.00238217f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.0405 $X2=0.7705 $Y2=0.0405
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7580 $Y=0.0405 $X2=0.7705 $Y2=0.0405
r3 9 5 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.7425
+ $Y=0.0405 $X2=0.7560 $Y2=0.0405
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.7275
+ $Y=0.0405 $X2=0.7425 $Y2=0.0405
r5 1 8 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.7020
+ $Y=0.0405 $X2=0.7275 $Y2=0.0405
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.0405 $X2=0.7000 $Y2=0.0405
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.0405 $X2=0.6875 $Y2=0.0405
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%SS VSS 9 31 40 12 10 11 4 15 3 14 1 16 13
c1 1 VSS 0.00106162f
c2 3 VSS 0.00610747f
c3 4 VSS 0.006775f
c4 9 VSS 0.0384426f
c5 10 VSS 0.00316024f
c6 11 VSS 0.00314802f
c7 12 VSS 0.0019167f
c8 13 VSS 0.0130321f
c9 14 VSS 0.00917009f
c10 15 VSS 0.0075344f
c11 16 VSS 0.00269071f
c12 17 VSS 0.00421859f
c13 18 VSS 0.00366088f
r1 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.2295 $X2=0.8620 $Y2=0.2295
r2 40 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.2295 $X2=0.8495 $Y2=0.2295
r3 4 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.2295
+ $X2=0.8640 $Y2=0.2340
r4 37 38 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.2340 $X2=0.8865 $Y2=0.2340
r5 14 18 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9180 $Y=0.2340 $X2=0.9450 $Y2=0.2340
r6 14 38 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.2340 $X2=0.8865 $Y2=0.2340
r7 18 35 6.74572 $w=1.545e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.2340 $X2=0.9450 $Y2=0.1980
r8 34 35 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1690 $X2=0.9450 $Y2=0.1980
r9 33 34 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1445 $X2=0.9450 $Y2=0.1690
r10 32 33 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1195 $X2=0.9450 $Y2=0.1445
r11 15 17 8.84443 $w=1.496e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.0810 $X2=0.9450 $Y2=0.0360
r12 15 32 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.0810 $X2=0.9450 $Y2=0.1195
r13 10 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.0405 $X2=0.8620 $Y2=0.0405
r14 31 10 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.0405 $X2=0.8495 $Y2=0.0405
r15 17 29 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.0360 $X2=0.9180 $Y2=0.0360
r16 3 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.0405
+ $X2=0.8640 $Y2=0.0360
r17 28 29 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.0360 $X2=0.9180 $Y2=0.0360
r18 27 28 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.0360 $X2=0.8910 $Y2=0.0360
r19 26 27 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.0360 $X2=0.8640 $Y2=0.0360
r20 13 16 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.0360 $X2=0.7830 $Y2=0.0360
r21 13 26 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0360 $X2=0.8370 $Y2=0.0360
r22 12 23 8.04505 $w=1.3e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.0705 $X2=0.7830 $Y2=0.1050
r23 12 16 6.39593 $w=1.55565e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7830 $Y=0.0705 $X2=0.7830 $Y2=0.0360
r24 1 20 2.36633 $w=2.3e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.7830
+ $Y=0.1055 $X2=0.7830 $Y2=0.1055
r25 1 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7830 $Y=0.1055
+ $X2=0.7830 $Y2=0.1050
r26 9 20 0.314665 $w=2.27e-07 $l=2.95e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.7830 $Y=0.1350 $X2=0.7830 $Y2=0.1055
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%MH VSS 9 47 51 57 61 10 3 16 20 1 17 4 12 14 18
+ 15 19
c1 1 VSS 0.000312446f
c2 3 VSS 0.00606346f
c3 4 VSS 0.00538477f
c4 9 VSS 0.036415f
c5 10 VSS 0.00226523f
c6 11 VSS 9.0832e-20
c7 12 VSS 0.00278446f
c8 13 VSS 6.982e-20
c9 14 VSS 0.00752837f
c10 15 VSS 0.00134331f
c11 16 VSS 0.000727687f
c12 17 VSS 0.000543512f
c13 18 VSS 0.00620285f
c14 19 VSS 2.27314e-20
c15 20 VSS 0.00279971f
r1 61 60 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r2 59 60 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r3 3 59 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3760 $Y=0.2295 $X2=0.3880 $Y2=0.2295
r4 13 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2295 $X2=0.3760 $Y2=0.2295
r5 55 56 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r6 57 55 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.1890 $X2=0.3635 $Y2=0.1890
r7 12 56 0.185185 $w=5.4e-08 $l=1e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r8 12 3 0.518519 $w=3.9e-08 $l=4.05494e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.1890 $X2=0.3760 $Y2=0.2295
r9 3 44 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2295
+ $X2=0.3780 $Y2=0.2340
r10 51 50 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r11 49 50 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4420 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r12 4 49 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4300 $Y=0.0405 $X2=0.4420 $Y2=0.0405
r13 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0405 $X2=0.4300 $Y2=0.0405
r14 10 4 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0810 $X2=0.4300 $Y2=0.0810
r15 47 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0810 $X2=0.4175 $Y2=0.0810
r16 44 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r17 42 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r18 41 42 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4160
+ $Y=0.2340 $X2=0.4050 $Y2=0.2340
r19 14 20 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4340
+ $Y=0.2340 $X2=0.4590 $Y2=0.2340
r20 14 41 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4340
+ $Y=0.2340 $X2=0.4160 $Y2=0.2340
r21 4 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0405
+ $X2=0.4320 $Y2=0.0360
r22 20 34 3.01468 $w=1.741e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4590 $Y2=0.2140
r23 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4455 $Y2=0.0360
r24 18 31 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4590 $Y2=0.0630
r25 18 37 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4455 $Y2=0.0360
r26 33 34 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1850 $X2=0.4590 $Y2=0.2140
r27 32 33 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1660 $X2=0.4590 $Y2=0.1850
r28 16 19 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1525 $X2=0.4590 $Y2=0.1310
r29 16 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1525 $X2=0.4590 $Y2=0.1660
r30 30 31 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0900 $X2=0.4590 $Y2=0.0630
r31 29 30 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1025 $X2=0.4590 $Y2=0.0900
r32 15 19 2.78392 $w=1.56471e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1140 $X2=0.4590 $Y2=0.1310
r33 15 29 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1140 $X2=0.4590 $Y2=0.1025
r34 19 27 4.18306 $w=1.49565e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1310 $X2=0.4820 $Y2=0.1310
r35 26 27 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5000
+ $Y=0.1310 $X2=0.4820 $Y2=0.1310
r36 25 26 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1310 $X2=0.5000 $Y2=0.1310
r37 17 24 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1310 $X2=0.5670 $Y2=0.1310
r38 17 25 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1310 $X2=0.5130 $Y2=0.1310
r39 23 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1330
+ $X2=0.5670 $Y2=0.1310
r40 1 22 1.47681 $w=1.53e-08 $l=9e-09 $layer=LIG $thickness=4.8e-08 $X=0.5670
+ $Y=0.1215 $X2=0.5670 $Y2=0.1305
r41 22 23 5.31651 $w=1.53e-08 $l=2.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.5670 $Y=0.1305 $X2=0.5670 $Y2=0.1330
r42 9 22 0.314665 $w=2.27e-07 $l=4.5e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5670 $Y=0.1350 $X2=0.5670 $Y2=0.1305
r43 3 12 1e-05
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%CLKN VSS 16 17 18 19 20 99 101 24 35 32 34 9 8
+ 22 21 26 25 1 27 36 23 29 2 5 30 10 3 28 31 33
c1 1 VSS 0.00146351f
c2 2 VSS 0.000295056f
c3 3 VSS 7.59612e-20
c4 4 VSS 1e-36
c5 5 VSS 0.000434637f
c6 8 VSS 0.00775466f
c7 9 VSS 0.0078539f
c8 10 VSS 0.00359183f
c9 16 VSS 0.0593859f
c10 17 VSS 0.00530001f
c11 18 VSS 0.00511876f
c12 19 VSS 0.00437364f
c13 20 VSS 0.00518215f
c14 21 VSS 0.00657876f
c15 22 VSS 0.00651999f
c16 23 VSS 0.00822253f
c17 24 VSS 0.00183535f
c18 25 VSS 0.00503549f
c19 26 VSS 0.00371036f
c20 27 VSS 0.000721628f
c21 28 VSS 0.000258222f
c22 29 VSS 0.000831314f
c23 30 VSS 0.00141386f
c24 31 VSS 0.00381093f
c25 32 VSS 0.00194944f
c26 33 VSS 0.00399733f
c27 34 VSS 0.000913807f
c28 35 VSS 0.000509073f
c29 36 VSS 0.0233792f
r1 101 100 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r2 22 100 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r3 99 98 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r4 21 98 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r5 9 96 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0550 $Y2=0.2340
r6 8 93 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0550 $Y2=0.0360
r7 95 96 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.2340 $X2=0.0550 $Y2=0.2340
r8 26 95 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0460 $Y2=0.2340
r9 26 33 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0180 $Y2=0.2340
r10 92 93 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.0360 $X2=0.0550 $Y2=0.0360
r11 25 92 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0460 $Y2=0.0360
r12 25 31 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0180 $Y2=0.0360
r13 5 91 2.78395 $w=2.4e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08 $X=0.7290
+ $Y=0.1780 $X2=0.7250 $Y2=0.1780
r14 20 5 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.7290 $Y=0.1350 $X2=0.7290 $Y2=0.1780
r15 4 84 10.3807 $w=2.30357e-08 $l=0 $layer=LISD $thickness=3.675e-08 $X=0.6210
+ $Y=0.1780 $X2=0.6210 $Y2=0.1780
r16 19 4 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.6210 $Y=0.1350 $X2=0.6210 $Y2=0.1780
r17 3 77 2.78395 $w=2.4e-08 $l=5e-09 $layer=LIG $thickness=4.8e-08 $X=0.4590
+ $Y=0.1780 $X2=0.4640 $Y2=0.1780
r18 18 3 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4590 $Y2=0.1780
r19 33 72 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.2340 $X2=0.0180 $Y2=0.2125
r20 31 71 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.0360 $X2=0.0180 $Y2=0.0575
r21 90 91 4.8113 $w=2.22e-08 $l=1.5e-09 $layer=LISD $thickness=2.7e-08
+ $X=0.7235 $Y=0.1780 $X2=0.7250 $Y2=0.1780
r22 89 90 10.8887 $w=2.22e-08 $l=2.15e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7020 $Y=0.1780 $X2=0.7235 $Y2=0.1780
r23 88 89 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6885 $Y=0.1780 $X2=0.7020 $Y2=0.1780
r24 87 88 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6750 $Y=0.1780 $X2=0.6885 $Y2=0.1780
r25 86 87 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6615 $Y=0.1780 $X2=0.6750 $Y2=0.1780
r26 85 86 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6480 $Y=0.1780 $X2=0.6615 $Y2=0.1780
r27 84 85 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6210 $Y=0.1780 $X2=0.6480 $Y2=0.1780
r28 83 84 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5940 $Y=0.1780 $X2=0.6210 $Y2=0.1780
r29 82 83 7.09034 $w=2.22e-08 $l=1.4e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5800 $Y=0.1780 $X2=0.5940 $Y2=0.1780
r30 81 82 6.58388 $w=2.22e-08 $l=1.3e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5670 $Y=0.1780 $X2=0.5800 $Y2=0.1780
r31 80 81 6.58388 $w=2.22e-08 $l=1.3e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5540 $Y=0.1780 $X2=0.5670 $Y2=0.1780
r32 79 80 7.09034 $w=2.22e-08 $l=1.4e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5400 $Y=0.1780 $X2=0.5540 $Y2=0.1780
r33 78 79 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5265 $Y=0.1780 $X2=0.5400 $Y2=0.1780
r34 76 77 10.3823 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4775 $Y=0.1780 $X2=0.4640 $Y2=0.1780
r35 75 76 11.142 $w=2.22e-08 $l=2.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4995 $Y=0.1780 $X2=0.4775 $Y2=0.1780
r36 74 78 1.51936 $w=2.22e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.5235
+ $Y=0.1780 $X2=0.5265 $Y2=0.1780
r37 73 74 5.31775 $w=2.22e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5130 $Y=0.1780 $X2=0.5235 $Y2=0.1780
r38 10 73 5.31775 $w=2.22e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5025 $Y=0.1780 $X2=0.5130 $Y2=0.1780
r39 10 75 1.51936 $w=2.22e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.5025
+ $Y=0.1780 $X2=0.4995 $Y2=0.1780
r40 2 65 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
r41 17 2 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r42 24 32 0.998523 $w=1.74118e-08 $l=1.01119e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1990 $X2=0.0165 $Y2=0.1890
r43 24 72 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1990 $X2=0.0180 $Y2=0.2125
r44 70 71 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0880 $X2=0.0180 $Y2=0.0575
r45 69 70 10.9599 $w=1.3e-08 $l=4.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1350 $X2=0.0180 $Y2=0.0880
r46 23 32 2.63085 $w=1.54194e-08 $l=1.7066e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1720 $X2=0.0165 $Y2=0.1890
r47 23 69 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1720 $X2=0.0180 $Y2=0.1350
r48 67 73 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5130 $Y=0.1845
+ $X2=0.5130 $Y2=0.1780
r49 30 67 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1680 $X2=0.5130 $Y2=0.1845
r50 65 66 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1555
r51 29 63 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1735 $X2=0.3510 $Y2=0.1890
r52 29 66 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1735 $X2=0.3510 $Y2=0.1555
r53 60 61 1.90199 $w=1.38333e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.0255 $Y=0.1890 $X2=0.0345 $Y2=0.1890
r54 32 60 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0165
+ $Y=0.1890 $X2=0.0255 $Y2=0.1890
r55 58 67 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.5130 $Y=0.1890
+ $X2=0.5130 $Y2=0.1845
r56 57 58 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.4320
+ $Y=0.1890 $X2=0.5130 $Y2=0.1890
r57 56 57 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1890 $X2=0.4320 $Y2=0.1890
r58 56 63 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.3510 $Y=0.1890
+ $X2=0.3510 $Y2=0.1890
r59 55 56 15.2739 $w=1.3e-08 $l=6.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.2855
+ $Y=0.1890 $X2=0.3510 $Y2=0.1890
r60 54 55 20.2875 $w=1.3e-08 $l=8.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.1985
+ $Y=0.1890 $X2=0.2855 $Y2=0.1890
r61 53 54 9.211 $w=1.3e-08 $l=3.95e-08 $layer=M2 $thickness=3.6e-08 $X=0.1590
+ $Y=0.1890 $X2=0.1985 $Y2=0.1890
r62 52 53 14.691 $w=1.3e-08 $l=6.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.0960
+ $Y=0.1890 $X2=0.1590 $Y2=0.1890
r63 51 52 14.691 $w=1.3e-08 $l=6.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.0330
+ $Y=0.1890 $X2=0.0960 $Y2=0.1890
r64 51 61 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.0330 $Y=0.1890
+ $X2=0.0345 $Y2=0.1890
r65 36 51 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.0215
+ $Y=0.1890 $X2=0.0330 $Y2=0.1890
r66 48 49 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1590
+ $Y=0.1890 $X2=0.1740 $Y2=0.1890
r67 48 53 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1590 $Y=0.1890
+ $X2=0.1590 $Y2=0.1890
r68 34 46 2.78392 $w=1.56471e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1890 $X2=0.1890 $Y2=0.1720
r69 34 49 2.31754 $w=1.6e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1890 $X2=0.1740 $Y2=0.1890
r70 28 35 2.78149 $w=1.76421e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1540 $X2=0.1890 $Y2=0.1350
r71 28 46 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1540 $X2=0.1890 $Y2=0.1720
r72 35 45 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1640 $Y2=0.1350
r73 44 45 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.1465
+ $Y=0.1350 $X2=0.1640 $Y2=0.1350
r74 43 44 0.46638 $w=1.3e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.1445
+ $Y=0.1350 $X2=0.1465 $Y2=0.1350
r75 42 43 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1445 $Y2=0.1350
r76 27 42 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1235
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r77 16 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r78 1 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
r79 9 22 1e-05
r80 8 21 1e-05
.ends

.subckt PM_DFFLQx4_ASAP7_75t_R%SH VSS 11 12 13 71 74 78 81 15 24 26 14 6 19 17
+ 18 5 16 22 2 28 27 21 23 1 25 20 29
c1 1 VSS 0.000693139f
c2 2 VSS 0.00780219f
c3 5 VSS 0.00473522f
c4 6 VSS 0.00527822f
c5 11 VSS 0.0374733f
c6 12 VSS 0.0810317f
c7 13 VSS 0.0809453f
c8 14 VSS 0.00498342f
c9 15 VSS 0.00516807f
c10 16 VSS 0.00788931f
c11 17 VSS 0.00193953f
c12 18 VSS 0.00190492f
c13 19 VSS 0.00262572f
c14 20 VSS 0.000823204f
c15 21 VSS 0.000471986f
c16 22 VSS 0.00133206f
c17 23 VSS 0.00261788f
c18 24 VSS 0.00688784f
c19 25 VSS 0.00270809f
c20 26 VSS 0.000154752f
c21 27 VSS 0.000399078f
c22 28 VSS 0.000378846f
c23 29 VSS 0.00981446f
r1 81 80 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r2 5 80 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6500 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r3 77 5 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6380 $Y=0.0405 $X2=0.6500 $Y2=0.0405
r4 14 77 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0405 $X2=0.6380 $Y2=0.0405
r5 78 14 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.0405 $X2=0.6335 $Y2=0.0405
r6 13 66 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=1.0530
+ $Y=0.1350 $X2=1.0530 $Y2=0.1360
r7 12 58 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.9990 $Y=0.1350 $X2=0.9990 $Y2=0.1360
r8 74 73 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r9 72 73 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7120 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r10 6 72 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7000 $Y=0.2295 $X2=0.7120 $Y2=0.2295
r11 15 6 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.2295 $X2=0.7000 $Y2=0.2295
r12 71 15 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.2295 $X2=0.6875 $Y2=0.2295
r13 5 56 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.0405
+ $X2=0.6480 $Y2=0.0360
r14 64 66 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.0405 $Y=0.1360 $X2=1.0530 $Y2=0.1360
r15 63 64 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.0260 $Y=0.1360 $X2=1.0405 $Y2=0.1360
r16 61 63 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.0115 $Y=0.1360 $X2=1.0260 $Y2=0.1360
r17 59 61 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=1.0085 $Y=0.1360 $X2=1.0115 $Y2=0.1360
r18 58 59 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.9990
+ $Y=0.1360 $X2=1.0085 $Y2=0.1360
r19 2 58 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.9895
+ $Y=0.1360 $X2=0.9990 $Y2=0.1360
r20 6 49 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7020 $Y=0.2295
+ $X2=0.7020 $Y2=0.2340
r21 56 57 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6480
+ $Y=0.0360 $X2=0.6615 $Y2=0.0360
r22 54 57 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0360 $X2=0.6615 $Y2=0.0360
r23 53 54 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6860
+ $Y=0.0360 $X2=0.6750 $Y2=0.0360
r24 16 25 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.7040
+ $Y=0.0360 $X2=0.7290 $Y2=0.0360
r25 16 53 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7040
+ $Y=0.0360 $X2=0.6860 $Y2=0.0360
r26 51 58 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.9990 $Y=0.1445
+ $X2=0.9990 $Y2=0.1360
r27 23 51 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.9990
+ $Y=0.1245 $X2=0.9990 $Y2=0.1445
r28 49 50 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.2340 $X2=0.7155 $Y2=0.2340
r29 24 50 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.2340 $X2=0.7155 $Y2=0.2340
r30 25 42 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.0360 $X2=0.7290 $Y2=0.0630
r31 46 51 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.9990 $Y=0.1530
+ $X2=0.9990 $Y2=0.1445
r32 45 46 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1530 $X2=0.9990 $Y2=0.1530
r33 44 45 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1530 $X2=0.9450 $Y2=0.1530
r34 29 44 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.8795
+ $Y=0.1530 $X2=0.8910 $Y2=0.1530
r35 43 44 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.8910 $Y=0.1485 $X2=0.8910
+ $Y2=0.1530
r36 22 43 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1305 $X2=0.8910 $Y2=0.1485
r37 18 38 6.50021 $w=1.33448e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1980 $X2=0.7290 $Y2=0.1690
r38 18 24 7.21452 $w=1.425e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1980 $X2=0.7290 $Y2=0.2340
r39 41 42 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.0900 $X2=0.7290 $Y2=0.0630
r40 40 41 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1090 $X2=0.7290 $Y2=0.0900
r41 17 26 4.67854 $w=1.44583e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1360 $X2=0.7290 $Y2=0.1600
r42 17 40 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1360 $X2=0.7290 $Y2=0.1090
r43 28 39 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1575 $X2=0.8910 $Y2=0.1665
r44 28 43 1.50855 $w=1.55e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1575 $X2=0.8910 $Y2=0.1485
r45 28 44 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.8910 $Y=0.1575 $X2=0.8910
+ $Y2=0.1530
r46 26 38 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1600 $X2=0.7290 $Y2=0.1690
r47 37 39 4.19024 $w=1.156e-08 $l=2.54018e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8660 $Y=0.1620 $X2=0.8910 $Y2=0.1665
r48 21 27 1.38478 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8480 $Y=0.1620 $X2=0.8370 $Y2=0.1620
r49 21 37 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8480
+ $Y=0.1620 $X2=0.8660 $Y2=0.1620
r50 36 38 4.4015 $w=1.35e-08 $l=2.78927e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7560 $Y=0.1620 $X2=0.7290 $Y2=0.1690
r51 35 36 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1620 $X2=0.7560 $Y2=0.1620
r52 19 27 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.1620 $X2=0.8370 $Y2=0.1620
r53 19 35 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.1620 $X2=0.7830 $Y2=0.1620
r54 27 34 4.88263 $w=1.47308e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8370 $Y=0.1620 $X2=0.8370 $Y2=0.1360
r55 20 34 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1180 $X2=0.8370 $Y2=0.1360
r56 33 34 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8370 $Y=0.1355
+ $X2=0.8370 $Y2=0.1360
r57 11 1 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.8370 $Y=0.1350 $X2=0.8370 $Y2=0.1245
r58 1 33 6.49795 $w=1.53e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08 $X=0.8370
+ $Y=0.1245 $X2=0.8370 $Y2=0.1355
.ends


*
.SUBCKT DFFLQx4_ASAP7_75t_R VSS VDD CLK D Q
*
* VSS VSS
* VDD VDD
* CLK CLK
* D D
* Q Q
*
*

MM20 N_MM20_d N_MM20_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM23 N_MM23_d N_MM22_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM10_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM6 N_MM6_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM12 N_MM12_d N_MM12_g N_MM12_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM17 N_MM17_d N_MM13_g N_MM17_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM16 N_MM16_d N_MM19_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM14 N_MM14_d N_MM14_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM24 N_MM24_d N_MM24_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@2 N_MM24@2_d N_MM24@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM0_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@4 N_MM0@4_d N_MM0@4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@3 N_MM0@3_d N_MM0@3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@2 N_MM0@2_d N_MM0@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM21 N_MM21_d N_MM20_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM22 N_MM22_d N_MM22_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM13 N_MM13_d N_MM13_g N_MM13_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM18 N_MM18_d N_MM18_g N_MM18_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM19 N_MM19_d N_MM19_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM15 N_MM15_d N_MM14_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM25 N_MM25_d N_MM24_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@2 N_MM25@2_d N_MM24@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2@4 N_MM2@4_d N_MM0@4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2@3 N_MM2@3_d N_MM0@3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2@2 N_MM2@2_d N_MM0@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "DFFLQx4_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "DFFLQx4_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_DFFLQx4_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_DFFLQx4_ASAP7_75t_R%noxref_24
cc_1 N_noxref_24_1 N_MM3_g 0.001371f
cc_2 N_noxref_24_1 N_CLKB_14 0.000770649f
cc_3 N_noxref_24_1 N_noxref_21_1 0.000470437f
cc_4 N_noxref_24_1 N_noxref_22_1 0.0077159f
cc_5 N_noxref_24_1 N_noxref_23_1 0.00123363f
x_PM_DFFLQx4_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_DFFLQx4_ASAP7_75t_R%noxref_23
cc_6 N_noxref_23_1 N_MM3_g 0.00136301f
cc_7 N_noxref_23_1 N_CLKB_13 0.000797653f
cc_8 N_noxref_23_1 N_noxref_21_1 0.00768789f
cc_9 N_noxref_23_1 N_noxref_22_1 0.000471705f
x_PM_DFFLQx4_ASAP7_75t_R%noxref_29 VSS N_noxref_29_1
+ PM_DFFLQx4_ASAP7_75t_R%noxref_29
cc_10 N_noxref_29_1 N_MM0@2_g 0.00146974f
cc_11 N_noxref_29_1 N_Q_14 0.000820809f
x_PM_DFFLQx4_ASAP7_75t_R%noxref_30 VSS N_noxref_30_1
+ PM_DFFLQx4_ASAP7_75t_R%noxref_30
cc_12 N_noxref_30_1 N_MM0@2_g 0.00147125f
cc_13 N_noxref_30_1 N_Q_16 0.000827762f
cc_14 N_noxref_30_1 N_noxref_29_1 0.00176533f
x_PM_DFFLQx4_ASAP7_75t_R%Q VSS Q N_MM0_d N_MM0@4_d N_MM0@3_d N_MM0@2_d
+ N_MM2@3_d N_MM2@2_d N_MM2_d N_MM2@4_d N_Q_14 N_Q_18 N_Q_16 N_Q_15 N_Q_13
+ N_Q_21 N_Q_20 N_Q_2 N_Q_3 N_Q_4 N_Q_1 PM_DFFLQx4_ASAP7_75t_R%Q
cc_15 N_Q_14 N_QN_1 0.000617754f
cc_16 N_Q_18 N_MM0@3_g 0.000637812f
cc_17 N_Q_16 N_MM0@3_g 0.0305264f
cc_18 N_Q_15 N_MM0_g 0.0306701f
cc_19 N_Q_13 N_MM0_g 0.0672379f
cc_20 N_Q_21 N_QN_22 0.00105722f
cc_21 N_Q_20 N_QN_20 0.00107359f
cc_22 N_Q_2 N_QN_19 0.00169079f
cc_23 N_Q_3 N_MM0@3_g 0.00183981f
cc_24 N_Q_4 N_MM0@3_g 0.00193267f
cc_25 N_Q_1 N_MM0_g 0.00222637f
cc_26 N_Q_2 N_MM0_g 0.00231359f
cc_27 N_Q_21 N_QN_18 0.00247263f
cc_28 N_Q_20 N_QN_17 0.00258346f
cc_29 N_Q_16 N_QN_1 0.00957989f
cc_30 N_Q_14 N_MM0@2_g 0.0367669f
cc_31 N_Q_13 N_MM0@4_g 0.0367911f
cc_32 N_Q_14 N_MM0@3_g 0.0700128f
x_PM_DFFLQx4_ASAP7_75t_R%noxref_28 VSS N_noxref_28_1
+ PM_DFFLQx4_ASAP7_75t_R%noxref_28
cc_33 N_noxref_28_1 N_SS_11 0.000654055f
cc_34 N_noxref_28_1 N_MM24_g 0.00171917f
cc_35 N_noxref_28_1 N_noxref_25_1 0.000477104f
cc_36 N_noxref_28_1 N_noxref_26_1 0.00776579f
cc_37 N_noxref_28_1 N_noxref_27_1 0.00123538f
x_PM_DFFLQx4_ASAP7_75t_R%noxref_26 VSS N_noxref_26_1
+ PM_DFFLQx4_ASAP7_75t_R%noxref_26
cc_38 N_noxref_26_1 N_SS_11 0.0169535f
cc_39 N_noxref_26_1 N_MM14_g 0.00619301f
cc_40 N_noxref_26_1 N_noxref_25_1 0.00153784f
x_PM_DFFLQx4_ASAP7_75t_R%QN VSS N_MM0_g N_MM0@4_g N_MM0@3_g N_MM0@2_g N_MM24_d
+ N_MM24@2_d N_MM25_d N_MM25@2_d N_QN_13 N_QN_16 N_QN_4 N_QN_17 N_QN_18 N_QN_14
+ N_QN_3 N_QN_1 N_QN_22 N_QN_20 N_QN_19 PM_DFFLQx4_ASAP7_75t_R%QN
cc_41 N_QN_13 N_SH_2 0.000391285f
cc_42 N_QN_13 N_SH_23 0.000639266f
cc_43 N_QN_13 N_MM24@2_g 0.0400009f
cc_44 N_QN_16 N_SH_23 0.000498905f
cc_45 N_QN_4 N_SH_2 0.000525096f
cc_46 N_QN_17 N_SH_2 0.000547453f
cc_47 N_QN_18 N_SH_2 0.000606613f
cc_48 N_QN_16 N_SH_29 0.000746558f
cc_49 N_QN_14 N_MM24_g 0.031445f
cc_50 N_QN_4 N_SH_23 0.00112025f
cc_51 N_MM0_g N_MM24@2_g 0.0016573f
cc_52 N_QN_3 N_MM24_g 0.0019584f
cc_53 N_QN_4 N_MM24_g 0.00211694f
cc_54 N_QN_14 N_SH_2 0.00514814f
cc_55 N_QN_13 N_MM24_g 0.069736f
x_PM_DFFLQx4_ASAP7_75t_R%noxref_27 VSS N_noxref_27_1
+ PM_DFFLQx4_ASAP7_75t_R%noxref_27
cc_56 N_noxref_27_1 N_SS_10 0.000649264f
cc_57 N_noxref_27_1 N_MM24_g 0.00171517f
cc_58 N_noxref_27_1 N_noxref_25_1 0.00777818f
cc_59 N_noxref_27_1 N_noxref_26_1 0.000482082f
x_PM_DFFLQx4_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_DFFLQx4_ASAP7_75t_R%noxref_25
cc_60 N_noxref_25_1 N_SS_10 0.0170443f
cc_61 N_noxref_25_1 N_MM14_g 0.00612547f
x_PM_DFFLQx4_ASAP7_75t_R%D VSS D N_MM3_g N_D_1 N_D_4 N_D_6 N_D_5
+ PM_DFFLQx4_ASAP7_75t_R%D
cc_62 N_MM3_g N_CLKN_29 0.000924367f
cc_63 N_D_1 N_CLKN_2 0.00230565f
cc_64 N_D_4 N_CLKN_36 0.000997757f
cc_65 N_D_4 N_CLKN_29 0.00436616f
cc_66 N_MM3_g N_MM1_g 0.00522658f
x_PM_DFFLQx4_ASAP7_75t_R%CLK VSS CLK N_MM20_g N_CLK_8 N_CLK_5 N_CLK_1 N_CLK_6
+ N_CLK_7 N_CLK_4 PM_DFFLQx4_ASAP7_75t_R%CLK
x_PM_DFFLQx4_ASAP7_75t_R%PD3 VSS N_MM9_s N_MM8_d N_PD3_1
+ PM_DFFLQx4_ASAP7_75t_R%PD3
cc_67 N_PD3_1 N_MM9_g 0.00776929f
cc_68 N_PD3_1 N_MM11_g 0.00769306f
x_PM_DFFLQx4_ASAP7_75t_R%PD2 VSS N_MM10_s N_MM11_d N_PD2_4 N_PD2_1 N_PD2_5
+ PM_DFFLQx4_ASAP7_75t_R%PD2
cc_69 N_PD2_4 N_CLKN_10 0.000148328f
cc_70 N_PD2_1 N_CLKN_3 0.000539312f
cc_71 N_PD2_5 N_CLKN_10 0.0012962f
cc_72 N_PD2_1 N_MM9_g 0.00208023f
cc_73 N_PD2_5 N_MM9_g 0.0073618f
cc_74 N_PD2_4 N_MM9_g 0.0239011f
cc_75 N_PD2_4 N_MM10_g 0.0149192f
cc_76 N_PD2_5 N_MM11_g 0.0147491f
cc_77 N_PD2_1 N_MH_16 0.00046468f
cc_78 N_PD2_4 N_MH_3 0.000601998f
cc_79 N_PD2_1 N_MH_20 0.00325091f
x_PM_DFFLQx4_ASAP7_75t_R%PU1 VSS N_MM3_d N_MM1_s N_PU1_1
+ PM_DFFLQx4_ASAP7_75t_R%PU1
cc_80 N_PU1_1 N_MM1_g 0.0169829f
cc_81 N_PU1_1 N_MM3_g 0.0172568f
x_PM_DFFLQx4_ASAP7_75t_R%PD4 VSS N_MM18_s N_MM19_d N_PD4_1
+ PM_DFFLQx4_ASAP7_75t_R%PD4
cc_82 N_PD4_1 N_MM18_g 0.00778436f
cc_83 N_PD4_1 N_MM19_g 0.00771036f
x_PM_DFFLQx4_ASAP7_75t_R%MS VSS N_MM11_g N_MM6_d N_MM12_d N_MM7_d N_MM13_d
+ N_MS_3 N_MS_15 N_MS_13 N_MS_12 N_MS_1 N_MS_17 N_MS_11 N_MS_4 N_MS_18 N_MS_14
+ N_MS_16 PM_DFFLQx4_ASAP7_75t_R%MS
cc_84 N_MS_3 N_CLKN_30 0.000222914f
cc_85 N_MS_3 N_CLKN_10 0.000582558f
cc_86 N_MS_3 N_CLKN_3 0.000126175f
cc_87 N_MS_3 N_MM9_g 0.000155367f
cc_88 N_MS_3 N_CLKN_36 0.000189619f
cc_89 N_MS_15 N_CLKN_30 0.000275548f
cc_90 N_MS_13 N_MM12_g 0.00788294f
cc_91 N_MS_12 N_MM12_g 0.00779054f
cc_92 N_MS_15 N_CLKN_10 0.000391047f
cc_93 N_MS_1 N_MM9_g 0.000568844f
cc_94 N_MS_17 N_CLKN_10 0.00155764f
cc_95 N_MS_11 N_MM12_g 0.00650573f
cc_96 N_MS_4 N_MM12_g 0.00257394f
cc_97 N_MS_4 N_CLKN_10 0.00631126f
cc_98 N_MM11_g N_MM9_g 0.0142133f
cc_99 N_MS_3 N_MM12_g 0.0259868f
cc_100 N_MS_13 N_MM10_g 0.000129f
cc_101 N_MS_13 N_CLKB_19 0.000367823f
cc_102 N_MS_13 N_CLKB_2 0.000210432f
cc_103 N_MS_13 N_CLKB_22 0.000242098f
cc_104 N_MS_17 N_CLKB_2 0.000265045f
cc_105 N_MS_17 N_CLKB_19 0.00443516f
cc_106 N_MS_18 N_CLKB_19 0.000663382f
cc_107 N_MS_14 N_CLKB_22 0.00267843f
cc_108 N_MS_13 N_MM13_g 0.0156027f
x_PM_DFFLQx4_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_DFFLQx4_ASAP7_75t_R%noxref_19
cc_109 N_noxref_19_1 N_MM20_g 0.00368134f
cc_110 N_noxref_19_1 N_CLKN_8 0.000541421f
cc_111 N_noxref_19_1 N_CLKN_9 4.19683e-20
cc_112 N_noxref_19_1 N_CLKN_31 5.93963e-20
cc_113 N_noxref_19_1 N_CLKN_23 0.000384397f
cc_114 N_noxref_19_1 N_CLKN_21 0.0276122f
x_PM_DFFLQx4_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_DFFLQx4_ASAP7_75t_R%noxref_21
cc_115 N_noxref_21_1 N_CLKN_1 0.000128874f
cc_116 N_noxref_21_1 N_MM22_g 0.00349545f
cc_117 N_noxref_21_1 N_CLKB_5 0.000442964f
cc_118 N_noxref_21_1 N_CLKB_13 0.0272531f
x_PM_DFFLQx4_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_DFFLQx4_ASAP7_75t_R%noxref_20
cc_119 N_noxref_20_1 N_MM20_g 0.00366879f
cc_120 N_noxref_20_1 N_CLKN_8 4.33592e-20
cc_121 N_noxref_20_1 N_CLKN_33 5.48613e-20
cc_122 N_noxref_20_1 N_CLKN_24 8.04419e-20
cc_123 N_noxref_20_1 N_CLKN_32 9.07629e-20
cc_124 N_noxref_20_1 N_CLKN_23 0.000271543f
cc_125 N_noxref_20_1 N_CLKN_9 0.000431355f
cc_126 N_noxref_20_1 N_CLKN_22 0.0275486f
cc_127 N_noxref_20_1 N_noxref_19_1 0.0020466f
x_PM_DFFLQx4_ASAP7_75t_R%PD1 VSS N_MM5_d N_MM4_s N_PD1_4 N_PD1_5 N_PD1_1
+ PM_DFFLQx4_ASAP7_75t_R%PD1
cc_128 N_PD1_4 N_CLKN_29 0.0002056f
cc_129 N_PD1_4 N_CLKN_2 0.00234205f
cc_130 N_PD1_4 N_MM1_g 0.0732719f
cc_131 N_PD1_4 N_D_1 0.000671945f
cc_132 N_PD1_4 N_D_4 0.000780487f
cc_133 N_PD1_4 N_MM3_g 0.0359455f
cc_134 N_PD1_5 N_CLKB_18 0.000307641f
cc_135 N_PD1_5 N_CLKB_1 0.000631522f
cc_136 N_PD1_5 N_MM10_g 0.0346046f
cc_137 N_PD1_1 N_MH_4 0.00121398f
cc_138 N_PD1_1 N_MH_10 0.00348095f
x_PM_DFFLQx4_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_DFFLQx4_ASAP7_75t_R%noxref_22
cc_139 N_noxref_22_1 N_CLKN_1 0.000125505f
cc_140 N_noxref_22_1 N_MM22_g 0.00363782f
cc_141 N_noxref_22_1 N_CLKB_6 0.000362156f
cc_142 N_noxref_22_1 N_CLKB_14 0.0271158f
cc_143 N_noxref_22_1 N_noxref_21_1 0.00146916f
x_PM_DFFLQx4_ASAP7_75t_R%CLKB VSS N_MM10_g N_MM13_g N_MM23_d N_MM22_d N_CLKB_17
+ N_CLKB_6 N_CLKB_5 N_CLKB_16 N_CLKB_15 N_CLKB_13 N_CLKB_21 N_CLKB_22 N_CLKB_14
+ N_CLKB_19 N_CLKB_18 N_CLKB_2 N_CLKB_1 N_CLKB_20 PM_DFFLQx4_ASAP7_75t_R%CLKB
cc_144 N_CLKB_17 N_CLK_5 9.56186e-20
cc_145 N_CLKB_6 N_CLK_5 0.000322611f
cc_146 N_CLKB_5 N_CLK_5 0.00043092f
cc_147 N_CLKB_16 N_CLK_5 0.000194943f
cc_148 N_CLKB_16 N_CLK_6 0.00096122f
cc_149 N_CLKB_15 N_CLK_5 0.0022788f
cc_150 N_CLKB_13 N_CLKN_25 3.79292e-20
cc_151 N_CLKB_13 N_CLKN_23 6.3854e-20
cc_152 N_MM13_g N_CLKN_5 0.000221483f
cc_153 N_CLKB_21 N_CLKN_34 0.000236989f
cc_154 N_CLKB_6 N_CLKN_34 0.000268926f
cc_155 N_CLKB_22 N_CLKN_30 0.000670286f
cc_156 N_CLKB_6 N_CLKN_1 0.000313272f
cc_157 N_CLKB_16 N_CLKN_34 0.00488981f
cc_158 N_CLKB_14 N_MM22_g 0.0111944f
cc_159 N_CLKB_15 N_CLKN_35 0.000459208f
cc_160 N_CLKB_22 N_CLKN_29 0.000528446f
cc_161 N_CLKB_19 N_CLKN_10 0.000550779f
cc_162 N_MM10_g N_CLKN_3 0.000562197f
cc_163 N_CLKB_18 N_CLKN_36 0.000609815f
cc_164 N_CLKB_14 N_CLKN_1 0.000622236f
cc_165 N_CLKB_2 N_CLKN_10 0.00268809f
cc_166 N_CLKB_6 N_CLKN_27 0.000715289f
cc_167 N_CLKB_5 N_MM22_g 0.000748735f
cc_168 N_CLKB_17 N_CLKN_36 0.000813788f
cc_169 N_CLKB_1 N_CLKN_2 0.00225507f
cc_170 N_CLKB_17 N_CLKN_28 0.000999347f
cc_171 N_CLKB_6 N_MM22_g 0.00110755f
cc_172 N_CLKB_18 N_CLKN_29 0.00313778f
cc_173 N_MM10_g N_MM9_g 0.0036824f
cc_174 N_CLKB_17 N_CLKN_35 0.0038056f
cc_175 N_MM13_g N_CLKN_10 0.00435676f
cc_176 N_MM13_g N_MM18_g 0.00583774f
cc_177 N_MM10_g N_MM1_g 0.00704712f
cc_178 N_MM13_g N_MM12_g 0.0182813f
cc_179 N_CLKB_22 N_CLKN_36 0.0280923f
cc_180 N_CLKB_13 N_MM22_g 0.0389085f
cc_181 N_CLKB_21 N_D_6 0.000702357f
cc_182 N_CLKB_20 N_D_5 0.00103036f
cc_183 N_CLKB_22 N_D_4 0.0011406f
cc_184 N_CLKB_17 N_D_4 0.00857312f
x_PM_DFFLQx4_ASAP7_75t_R%PD5 VSS N_MM17_s N_MM16_d N_PD5_1 N_PD5_5 N_PD5_4
+ PM_DFFLQx4_ASAP7_75t_R%PD5
cc_185 N_PD5_1 N_MM18_g 0.000854635f
cc_186 N_PD5_5 N_MM18_g 0.00694921f
cc_187 N_PD5_4 N_MM18_g 0.0240453f
cc_188 N_PD5_4 N_MM13_g 0.0153104f
cc_189 N_PD5_1 N_MM19_g 0.000898764f
cc_190 N_PD5_5 N_MM19_g 0.0156146f
cc_191 N_PD5_1 N_SH_14 0.000317886f
cc_192 N_PD5_1 N_SH_16 0.000455708f
cc_193 N_PD5_1 N_SH_17 0.000564907f
cc_194 N_PD5_4 N_SH_5 0.000657708f
cc_195 N_PD5_1 N_SH_25 0.00253443f
x_PM_DFFLQx4_ASAP7_75t_R%SS VSS N_MM19_g N_MM14_d N_MM15_d N_SS_12 N_SS_10
+ N_SS_11 N_SS_4 N_SS_15 N_SS_3 N_SS_14 N_SS_1 N_SS_16 N_SS_13
+ PM_DFFLQx4_ASAP7_75t_R%SS
cc_196 N_MM19_g N_CLKN_10 0.000223052f
cc_197 N_MM19_g N_CLKN_5 0.000532379f
cc_198 N_MM19_g N_MM18_g 0.0135188f
x_PM_DFFLQx4_ASAP7_75t_R%MH VSS N_MM7_g N_MM4_d N_MM9_d N_MM1_d N_MM10_d
+ N_MH_10 N_MH_3 N_MH_16 N_MH_20 N_MH_1 N_MH_17 N_MH_4 N_MH_12 N_MH_14 N_MH_18
+ N_MH_15 N_MH_19 PM_DFFLQx4_ASAP7_75t_R%MH
cc_199 N_MH_10 N_CLKN_30 0.000392195f
cc_200 N_MH_10 N_MM1_g 0.000431834f
cc_201 N_MH_10 N_CLKN_29 0.000370343f
cc_202 N_MH_3 N_CLKN_2 0.000279932f
cc_203 N_MH_16 N_CLKN_30 0.00277617f
cc_204 N_MH_20 N_CLKN_30 0.000312674f
cc_205 N_MH_1 N_CLKN_10 0.00211017f
cc_206 N_MH_17 N_CLKN_10 0.000621675f
cc_207 N_MH_4 N_MM9_g 0.000634053f
cc_208 N_MH_12 N_CLKN_2 0.000787943f
cc_209 N_MH_16 N_CLKN_3 0.000792291f
cc_210 N_MH_3 N_CLKN_29 0.00138981f
cc_211 N_MH_14 N_CLKN_29 0.00141058f
cc_212 N_MH_14 N_CLKN_36 0.00151164f
cc_213 N_MH_3 N_MM1_g 0.00177427f
cc_214 N_MH_17 N_CLKN_30 0.00362455f
cc_215 N_MM7_g N_CLKN_10 0.00460892f
cc_216 N_MH_12 N_MM1_g 0.0336855f
cc_217 N_MM7_g N_MM12_g 0.0127547f
cc_218 N_MH_10 N_MM9_g 0.0363712f
cc_219 N_MH_10 N_CLKB_2 0.000100568f
cc_220 N_MH_10 N_MM13_g 0.000161062f
cc_221 N_MH_10 N_CLKB_18 0.000273899f
cc_222 N_MH_14 N_CLKB_18 0.000341422f
cc_223 N_MH_18 N_CLKB_18 0.000363029f
cc_224 N_MH_12 N_MM10_g 0.0163831f
cc_225 N_MH_3 N_CLKB_1 0.000825608f
cc_226 N_MH_4 N_MM10_g 0.00108808f
cc_227 N_MH_15 N_CLKB_18 0.00116335f
cc_228 N_MH_3 N_MM10_g 0.00117127f
cc_229 N_MH_17 N_CLKB_22 0.0012439f
cc_230 N_MH_16 N_CLKB_18 0.00127122f
cc_231 N_MH_12 N_CLKB_1 0.00160994f
cc_232 N_MH_16 N_CLKB_22 0.00230808f
cc_233 N_MH_19 N_CLKB_18 0.0028802f
cc_234 N_MH_10 N_MM10_g 0.053063f
cc_235 N_MH_4 N_MS_1 0.000402005f
cc_236 N_MH_17 N_MS_18 0.000564066f
cc_237 N_MH_17 N_MS_1 0.000817588f
cc_238 N_MM7_g N_MS_3 0.000981901f
cc_239 N_MH_17 N_MS_17 0.00100661f
cc_240 N_MH_1 N_MS_14 0.00104006f
cc_241 N_MH_1 N_MM11_g 0.00107124f
cc_242 N_MM7_g N_MS_1 0.00116091f
cc_243 N_MH_15 N_MS_14 0.00126889f
cc_244 N_MM7_g N_MS_12 0.00633515f
cc_245 N_MM7_g N_MS_11 0.00641993f
cc_246 N_MH_17 N_MS_14 0.00715447f
cc_247 N_MM7_g N_MM11_g 0.02949f
x_PM_DFFLQx4_ASAP7_75t_R%CLKN VSS N_MM22_g N_MM1_g N_MM9_g N_MM12_g N_MM18_g
+ N_MM20_d N_MM21_d N_CLKN_24 N_CLKN_35 N_CLKN_32 N_CLKN_34 N_CLKN_9 N_CLKN_8
+ N_CLKN_22 N_CLKN_21 N_CLKN_26 N_CLKN_25 N_CLKN_1 N_CLKN_27 N_CLKN_36
+ N_CLKN_23 N_CLKN_29 N_CLKN_2 N_CLKN_5 N_CLKN_30 N_CLKN_10 N_CLKN_3 N_CLKN_28
+ N_CLKN_31 N_CLKN_33 PM_DFFLQx4_ASAP7_75t_R%CLKN
cc_248 N_CLKN_24 N_MM20_g 7.87466e-20
cc_249 N_CLKN_35 N_MM20_g 8.63073e-20
cc_250 N_CLKN_32 N_MM20_g 0.000193835f
cc_251 N_CLKN_34 N_MM20_g 0.000204278f
cc_252 N_CLKN_9 N_MM20_g 0.00111872f
cc_253 N_CLKN_8 N_MM20_g 0.00117142f
cc_254 N_CLKN_22 N_MM20_g 0.0112145f
cc_255 N_CLKN_21 N_MM20_g 0.0112238f
cc_256 N_CLKN_26 N_CLK_8 0.000654695f
cc_257 N_CLKN_25 N_CLK_5 0.000782923f
cc_258 N_CLKN_1 N_CLK_8 0.000904332f
cc_259 N_CLKN_27 N_CLK_1 0.000916011f
cc_260 N_CLKN_26 N_CLK_6 0.00130298f
cc_261 N_CLKN_27 N_CLK_7 0.00139414f
cc_262 N_CLKN_36 N_CLK_8 0.00170362f
cc_263 N_CLKN_23 N_CLK_4 0.00176918f
cc_264 N_CLKN_27 N_CLK_4 0.00200673f
cc_265 N_CLKN_34 N_CLK_8 0.00228058f
cc_266 N_CLKN_1 N_CLK_1 0.0023354f
cc_267 N_CLKN_25 N_CLK_7 0.00234697f
cc_268 N_CLKN_27 N_CLK_8 0.00247431f
cc_269 N_CLKN_32 N_CLK_8 0.00259441f
cc_270 N_MM22_g N_MM20_g 0.0351335f
x_PM_DFFLQx4_ASAP7_75t_R%SH VSS N_MM14_g N_MM24_g N_MM24@2_g N_MM13_s N_MM18_d
+ N_MM12_s N_MM17_d N_SH_15 N_SH_24 N_SH_26 N_SH_14 N_SH_6 N_SH_19 N_SH_17
+ N_SH_18 N_SH_5 N_SH_16 N_SH_22 N_SH_2 N_SH_28 N_SH_27 N_SH_21 N_SH_23 N_SH_1
+ N_SH_25 N_SH_20 N_SH_29 PM_DFFLQx4_ASAP7_75t_R%SH
cc_271 N_SH_15 N_CLKN_36 0.000102705f
cc_272 N_SH_24 N_CLKN_10 0.000172976f
cc_273 N_SH_26 N_CLKN_10 0.000209498f
cc_274 N_SH_14 N_MM12_g 0.00680269f
cc_275 N_SH_6 N_CLKN_10 0.000290006f
cc_276 N_SH_19 N_CLKN_5 0.000420754f
cc_277 N_SH_17 N_CLKN_10 0.000427359f
cc_278 N_SH_18 N_CLKN_10 0.00058065f
cc_279 N_SH_15 N_CLKN_5 0.000925729f
cc_280 N_SH_6 N_MM18_g 0.00098771f
cc_281 N_SH_15 N_CLKN_10 0.00224933f
cc_282 N_SH_5 N_MM12_g 0.00950874f
cc_283 N_SH_15 N_MM18_g 0.0161875f
cc_284 N_SH_5 N_CLKB_22 0.000127335f
cc_285 N_SH_6 N_MM13_g 0.000165609f
cc_286 N_SH_19 N_CLKB_19 0.00021532f
cc_287 N_SH_14 N_MM13_g 0.00677f
cc_288 N_SH_15 N_MM13_g 0.00683705f
cc_289 N_SH_24 N_CLKB_19 0.00032371f
cc_290 N_SH_26 N_CLKB_19 0.000945636f
cc_291 N_SH_17 N_CLKB_2 0.000447194f
cc_292 N_SH_18 N_CLKB_19 0.000527203f
cc_293 N_SH_5 N_CLKB_2 0.000527576f
cc_294 N_SH_16 N_CLKB_19 0.000527852f
cc_295 N_SH_16 N_CLKB_22 0.00106945f
cc_296 N_SH_17 N_CLKB_19 0.00400914f
cc_297 N_SH_5 N_MM13_g 0.0184242f
cc_298 N_SH_17 N_MS_3 0.000113584f
cc_299 N_SH_24 N_MS_3 0.000157802f
cc_300 N_SH_15 N_MS_3 0.00043608f
cc_301 N_SH_14 N_MS_3 0.000466061f
cc_302 N_SH_6 N_MS_3 0.000247552f
cc_303 N_SH_24 N_MS_4 0.000292847f
cc_304 N_SH_6 N_MS_4 0.000422215f
cc_305 N_SH_24 N_MS_17 0.00054474f
cc_306 N_SH_15 N_MS_4 0.000586083f
cc_307 N_SH_16 N_MS_16 0.000589783f
cc_308 N_SH_16 N_MS_18 0.00161483f
cc_309 N_SH_5 N_MS_3 0.00367235f
cc_310 N_SH_18 N_MM19_g 0.000145864f
cc_311 N_SH_22 N_MM19_g 0.000149903f
cc_312 N_SH_2 N_MM19_g 0.000157237f
cc_313 N_SH_28 N_MM19_g 0.000158627f
cc_314 N_SH_27 N_SS_12 0.000212455f
cc_315 N_MM14_g N_SS_10 0.00676597f
cc_316 N_MM14_g N_SS_11 0.00687672f
cc_317 N_SH_21 N_SS_4 0.000262972f
cc_318 N_SH_2 N_SS_15 0.000282312f
cc_319 N_SH_23 N_SS_15 0.00154401f
cc_320 N_SH_22 N_SS_15 0.00674405f
cc_321 N_MM14_g N_SS_3 0.000400856f
cc_322 N_MM14_g N_SS_4 0.000514006f
cc_323 N_SH_21 N_SS_14 0.000659397f
cc_324 N_SH_1 N_SS_1 0.000700509f
cc_325 N_SH_25 N_SS_16 0.000833035f
cc_326 N_SH_17 N_SS_1 0.000845703f
cc_327 N_SH_28 N_SS_15 0.000909051f
cc_328 N_SH_20 N_SS_12 0.000981574f
cc_329 N_SH_20 N_SS_13 0.000994696f
cc_330 N_MM14_g N_SS_1 0.00110489f
cc_331 N_SH_1 N_MM19_g 0.00113976f
cc_332 N_SH_28 N_SS_14 0.00133107f
cc_333 N_SH_19 N_SS_12 0.00157373f
cc_334 N_SH_29 N_SS_15 0.00187294f
cc_335 N_SH_17 N_SS_12 0.00489906f
cc_336 N_MM14_g N_MM19_g 0.0294844f
*END of DFFLQx4_ASAP7_75t_R.pxi
.ENDS
** Design:	SDFHx1_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "SDFHx1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "SDFHx1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_SDFHx1_ASAP7_75t_R%NET0166 VSS 2 3 1
c1 1 VSS 0.000995403f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3780 $Y2=0.0675
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%noxref_31 VSS 1
c1 1 VSS 0.00358062f
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%noxref_32 VSS 1
c1 1 VSS 0.00379131f
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%noxref_33 VSS 1
c1 1 VSS 0.00358767f
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%noxref_34 VSS 1
c1 1 VSS 0.00397078f
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%NET0167 VSS 14 28 7 9 1 11 12 10 8 2
c1 1 VSS 0.00638701f
c2 2 VSS 0.00553597f
c3 7 VSS 0.00465831f
c4 8 VSS 0.00319625f
c5 9 VSS 0.000965946f
c6 10 VSS 0.0175163f
c7 11 VSS 0.00163471f
c8 12 VSS 0.00204199f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0675 $X2=0.4840 $Y2=0.0675
r2 28 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4715 $Y2=0.0675
r3 2 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0675
+ $X2=0.4860 $Y2=0.0360
r4 24 25 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4475
+ $Y=0.0360 $X2=0.4860 $Y2=0.0360
r5 23 24 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4160
+ $Y=0.0360 $X2=0.4475 $Y2=0.0360
r6 22 23 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0360 $X2=0.4160 $Y2=0.0360
r7 21 22 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.3875
+ $Y=0.0360 $X2=0.4050 $Y2=0.0360
r8 20 21 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3605
+ $Y=0.0360 $X2=0.3875 $Y2=0.0360
r9 19 20 7.92845 $w=1.3e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3265
+ $Y=0.0360 $X2=0.3605 $Y2=0.0360
r10 10 12 1.03257 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3085 $Y=0.0360 $X2=0.2970 $Y2=0.0360
r11 10 19 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3085
+ $Y=0.0360 $X2=0.3265 $Y2=0.0360
r12 12 18 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.2970 $Y2=0.0540
r13 9 17 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0720 $X2=0.2970 $Y2=0.0900
r14 9 18 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0720 $X2=0.2970 $Y2=0.0540
r15 16 17 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2835 $Y=0.0900 $X2=0.2970 $Y2=0.0900
r16 11 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0900 $X2=0.2835 $Y2=0.0900
r17 11 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0900
+ $X2=0.2700 $Y2=0.0945
r18 1 15 23.8708 $w=2.02e-08 $l=4.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.2700 $Y=0.0540 $X2=0.2700 $Y2=0.0945
r19 14 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r20 7 13 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r21 1 7 1e-05
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%noxref_35 VSS 1
c1 1 VSS 0.00468338f
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%noxref_36 VSS 1
c1 1 VSS 0.00459056f
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%QN VSS 19 13 25 10 7 11 2 1 8 9
c1 1 VSS 0.00819579f
c2 2 VSS 0.00824718f
c3 7 VSS 0.00366303f
c4 8 VSS 0.00364396f
c5 9 VSS 0.00327762f
c6 10 VSS 0.00557949f
c7 11 VSS 0.00633277f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.2815 $Y=0.2025 $X2=1.2940 $Y2=0.2025
r2 25 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.2790 $Y=0.2025 $X2=1.2815 $Y2=0.2025
r3 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.2960 $Y=0.2025
+ $X2=1.2960 $Y2=0.2340
r4 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.2960
+ $Y=0.2340 $X2=1.3095 $Y2=0.2340
r5 11 20 1.09329 $w=1.76154e-08 $l=9.8e-09 $layer=M1 $thickness=3.6e-08
+ $X=1.3230 $Y=0.2340 $X2=1.3230 $Y2=0.2242
r6 11 23 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3230 $Y=0.2340 $X2=1.3095 $Y2=0.2340
r7 19 20 0.291487 $w=1.3e-08 $l=1.2e-09 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.2230 $X2=1.3230 $Y2=0.2242
r8 19 18 2.73998 $w=1.3e-08 $l=1.18e-08 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.2230 $X2=1.3230 $Y2=0.2112
r9 17 18 15.4488 $w=1.3e-08 $l=6.62e-08 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.1450 $X2=1.3230 $Y2=0.2112
r10 9 16 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3230 $Y=0.0675 $X2=1.3230 $Y2=0.0360
r11 9 17 18.0722 $w=1.3e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.0675 $X2=1.3230 $Y2=0.1450
r12 15 16 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3095 $Y=0.0360 $X2=1.3230 $Y2=0.0360
r13 14 15 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.2960
+ $Y=0.0360 $X2=1.3095 $Y2=0.0360
r14 10 14 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.2845
+ $Y=0.0360 $X2=1.2960 $Y2=0.0360
r15 1 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.2960 $Y=0.0675
+ $X2=1.2960 $Y2=0.0360
r16 7 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.2815 $Y=0.0675 $X2=1.2940 $Y2=0.0675
r17 13 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.2790 $Y=0.0675 $X2=1.2815 $Y2=0.0675
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.00425088f
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.00434087f
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%D VSS 11 3 5 4 1
c1 1 VSS 0.00675184f
c2 3 VSS 0.0458469f
c3 4 VSS 0.005878f
c4 5 VSS 0.00442473f
r1 11 5 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M2 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1170 $X2=0.3665 $Y2=0.1170
r2 11 9 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4050 $Y=0.1170 $X2=0.4050
+ $Y2=0.1170
r3 4 9 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1170
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r5 1 4 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%SEN VSS 9 48 50 16 12 14 4 10 11 13 3 1 15
c1 1 VSS 0.00389808f
c2 3 VSS 0.00854277f
c3 4 VSS 0.00686379f
c4 9 VSS 0.0815442f
c5 10 VSS 0.00425337f
c6 11 VSS 0.00458575f
c7 12 VSS 0.00170371f
c8 13 VSS 0.00372935f
c9 14 VSS 0.000832184f
c10 15 VSS 0.00589979f
c11 16 VSS 0.0132551f
r1 50 49 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.2050 $Y=0.2295 $X2=1.2025 $Y2=0.2295
r2 11 49 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.1900 $Y=0.2295 $X2=1.2025 $Y2=0.2295
r3 4 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.1880 $Y=0.2295
+ $X2=1.1880 $Y2=0.2340
r4 48 47 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.2050 $Y=0.0405 $X2=1.2025 $Y2=0.0405
r5 10 47 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.1900 $Y=0.0405 $X2=1.2025 $Y2=0.0405
r6 44 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.1745
+ $Y=0.2340 $X2=1.1880 $Y2=0.2340
r7 15 40 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1610 $Y=0.2340 $X2=1.1610 $Y2=0.2125
r8 15 44 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1610 $Y=0.2340 $X2=1.1745 $Y2=0.2340
r9 42 10 3.98201 $w=3.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.1730 $Y=0.0455 $X2=1.1880 $Y2=0.0455
r10 41 42 3.18561 $w=3.32e-08 $l=1.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.1610 $Y=0.0455 $X2=1.1730 $Y2=0.0455
r11 3 41 3.31834 $w=3.32e-08 $l=1.25e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.1485 $Y=0.0455 $X2=1.1610 $Y2=0.0455
r12 39 40 15.7403 $w=1.3e-08 $l=6.75e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.1450 $X2=1.1610 $Y2=0.2125
r13 38 39 14.9241 $w=1.3e-08 $l=6.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0810 $X2=1.1610 $Y2=0.1450
r14 37 38 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0650 $X2=1.1610 $Y2=0.0810
r15 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0515 $X2=1.1610 $Y2=0.0650
r16 36 41 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.1610 $Y=0.0515
+ $X2=1.1610 $Y2=0.0455
r17 35 36 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0425 $X2=1.1610 $Y2=0.0515
r18 13 35 1.28254 $w=1.3e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0370 $X2=1.1610 $Y2=0.0425
r19 33 38 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=1.1610 $Y=0.0810
+ $X2=1.1610 $Y2=0.0810
r20 32 33 27.2832 $w=1.3e-08 $l=1.17e-07 $layer=M2 $thickness=3.6e-08 $X=1.0440
+ $Y=0.0810 $X2=1.1610 $Y2=0.0810
r21 31 32 29.3819 $w=1.3e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.9180
+ $Y=0.0810 $X2=1.0440 $Y2=0.0810
r22 30 31 40.3418 $w=1.3e-08 $l=1.73e-07 $layer=M2 $thickness=3.6e-08 $X=0.7450
+ $Y=0.0810 $X2=0.9180 $Y2=0.0810
r23 29 30 50.4856 $w=1.3e-08 $l=2.165e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.5285 $Y=0.0810 $X2=0.7450 $Y2=0.0810
r24 28 29 17.9556 $w=1.3e-08 $l=7.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.4515
+ $Y=0.0810 $X2=0.5285 $Y2=0.0810
r25 27 28 12.4757 $w=1.3e-08 $l=5.35e-08 $layer=M2 $thickness=3.6e-08 $X=0.3980
+ $Y=0.0810 $X2=0.4515 $Y2=0.0810
r26 26 27 10.9599 $w=1.3e-08 $l=4.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0810 $X2=0.3980 $Y2=0.0810
r27 16 26 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.3395
+ $Y=0.0810 $X2=0.3510 $Y2=0.0810
r28 14 22 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.0720 $X2=0.3510 $Y2=0.0855
r29 14 26 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.3510 $Y=0.0720 $X2=0.3510
+ $Y2=0.0810
r30 22 23 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0855 $X2=0.3510 $Y2=0.0945
r31 22 26 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.3510 $Y=0.0855 $X2=0.3510
+ $Y2=0.0810
r32 21 23 1.86552 $w=1.3e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1025 $X2=0.3510 $Y2=0.0945
r33 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1160 $X2=0.3510 $Y2=0.1025
r34 12 20 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1160
r35 9 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r36 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
r37 4 11 1e-05
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%CLK VSS 14 3 6 8 1 5 4 7
c1 1 VSS 0.00260449f
c2 3 VSS 0.0597449f
c3 4 VSS 0.00123214f
c4 5 VSS 0.00457896f
c5 6 VSS 0.00167991f
c6 7 VSS 0.00126307f
c7 8 VSS 0.00437414f
r1 8 18 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.1940 $X2=0.0945 $Y2=0.1940
r2 5 17 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0630 $X2=0.1080 $Y2=0.0900
r3 7 15 1.44308 $w=1.7e-08 $l=1.13e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1940 $X2=0.0810 $Y2=0.1827
r4 7 18 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1940 $X2=0.0945 $Y2=0.1940
r5 16 17 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.0900 $X2=0.1080 $Y2=0.0900
r6 6 16 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0900 $X2=0.0945 $Y2=0.0900
r7 14 15 0.641272 $w=1.3e-08 $l=2.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1800 $X2=0.0810 $Y2=0.1827
r8 14 13 1.57403 $w=1.3e-08 $l=6.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1800 $X2=0.0810 $Y2=0.1732
r9 12 13 4.13912 $w=1.3e-08 $l=1.77e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1555 $X2=0.0810 $Y2=0.1732
r10 11 12 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1555
r11 10 11 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1235 $X2=0.0810 $Y2=0.1350
r12 4 10 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1100 $X2=0.0810 $Y2=0.1235
r13 4 6 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1100 $X2=0.0810 $Y2=0.0900
r14 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r15 1 11 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%NET0141 VSS 12 13 27 28 7 9 1 8 2
c1 1 VSS 0.00531812f
c2 2 VSS 0.00527243f
c3 7 VSS 0.003341f
c4 8 VSS 0.00337113f
c5 9 VSS 0.00264182f
r1 28 26 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r2 2 26 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r4 27 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r5 2 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.1980
r6 22 23 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4205
+ $Y=0.1980 $X2=0.4320 $Y2=0.1980
r7 21 22 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4160
+ $Y=0.1980 $X2=0.4205 $Y2=0.1980
r8 20 21 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1980 $X2=0.4160 $Y2=0.1980
r9 19 20 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.3875
+ $Y=0.1980 $X2=0.4050 $Y2=0.1980
r10 18 19 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3695
+ $Y=0.1980 $X2=0.3875 $Y2=0.1980
r11 17 18 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1980 $X2=0.3695 $Y2=0.1980
r12 16 17 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.1980 $X2=0.3510 $Y2=0.1980
r13 15 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1980 $X2=0.3375 $Y2=0.1980
r14 14 15 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3130
+ $Y=0.1980 $X2=0.3240 $Y2=0.1980
r15 9 14 0.699569 $w=1.3e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.3100
+ $Y=0.1980 $X2=0.3130 $Y2=0.1980
r16 1 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.1980
r17 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r18 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r19 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r20 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%CLKN VSS 13 14 15 71 73 8 18 7 17 16 19 1 23 25
+ 22 21 20 3 2 24
c1 1 VSS 0.00139529f
c2 2 VSS 0.000108846f
c3 3 VSS 0.000191667f
c4 7 VSS 0.00789574f
c5 8 VSS 0.00784343f
c6 13 VSS 0.059311f
c7 14 VSS 0.00448367f
c8 15 VSS 0.00460295f
c9 16 VSS 0.006288f
c10 17 VSS 0.00620181f
c11 18 VSS 0.0106232f
c12 19 VSS 0.000480532f
c13 20 VSS 0.000101498f
c14 21 VSS 0.00048105f
c15 22 VSS 0.00779123f
c16 23 VSS 0.00672242f
c17 24 VSS 0.000163452f
c18 25 VSS 0.0209278f
r1 73 72 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r2 17 72 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r3 71 70 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r4 16 70 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r5 8 66 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0540 $Y2=0.2340
r6 7 63 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0540 $Y2=0.0360
r7 1 58 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1440
r8 13 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r9 65 66 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r10 23 57 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.2340 $X2=0.0270 $Y2=0.2140
r11 23 65 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0405 $Y2=0.2340
r12 62 63 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r13 22 55 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0360 $X2=0.0270 $Y2=0.0630
r14 22 62 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0360 $X2=0.0405 $Y2=0.0360
r15 2 49 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6210 $Y=0.1350
+ $X2=0.6210 $Y2=0.1395
r16 14 2 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1350
r17 19 58 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1235 $X2=0.1350 $Y2=0.1440
r18 56 57 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1940 $X2=0.0270 $Y2=0.2140
r19 54 55 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0900 $X2=0.0270 $Y2=0.0630
r20 53 56 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1735 $X2=0.0270 $Y2=0.1940
r21 52 53 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1530 $X2=0.0270 $Y2=0.1735
r22 18 52 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1215 $X2=0.0270 $Y2=0.1530
r23 18 54 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1215 $X2=0.0270 $Y2=0.0900
r24 24 49 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1620 $X2=0.6210 $Y2=0.1395
r25 24 37 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.6210 $Y=0.1620 $X2=0.6210
+ $Y2=0.1530
r26 20 49 5.47996 $w=1.3e-08 $l=2.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1160 $X2=0.6210 $Y2=0.1395
r27 47 48 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1530 $X2=0.1595 $Y2=0.1530
r28 47 58 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1350 $Y=0.1530
+ $X2=0.1350 $Y2=0.1440
r29 46 47 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1530 $X2=0.1350 $Y2=0.1530
r30 45 46 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1530 $X2=0.0810 $Y2=0.1530
r31 45 52 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.0270 $Y=0.1530
+ $X2=0.0270 $Y2=0.1530
r32 43 48 7.81186 $w=1.3e-08 $l=3.35e-08 $layer=M2 $thickness=3.6e-08 $X=0.1930
+ $Y=0.1530 $X2=0.1595 $Y2=0.1530
r33 42 43 12.7088 $w=1.3e-08 $l=5.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.2475
+ $Y=0.1530 $X2=0.1930 $Y2=0.1530
r34 41 42 26.2338 $w=1.3e-08 $l=1.125e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.3600 $Y=0.1530 $X2=0.2475 $Y2=0.1530
r35 40 41 21.3369 $w=1.3e-08 $l=9.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.4515
+ $Y=0.1530 $X2=0.3600 $Y2=0.1530
r36 39 40 17.9556 $w=1.3e-08 $l=7.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.5285
+ $Y=0.1530 $X2=0.4515 $Y2=0.1530
r37 37 38 15.2739 $w=1.3e-08 $l=6.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1530 $X2=0.6865 $Y2=0.1530
r38 37 49 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.6210 $Y=0.1530 $X2=0.6210
+ $Y2=0.1395
r39 36 37 4.6638 $w=1.3e-08 $l=2e-08 $layer=M2 $thickness=3.6e-08 $X=0.6010
+ $Y=0.1530 $X2=0.6210 $Y2=0.1530
r40 36 39 16.9063 $w=1.3e-08 $l=7.25e-08 $layer=M2 $thickness=3.6e-08 $X=0.6010
+ $Y=0.1530 $X2=0.5285 $Y2=0.1530
r41 25 35 18.3054 $w=1.3e-08 $l=7.85e-08 $layer=M2 $thickness=3.6e-08 $X=0.8125
+ $Y=0.1530 $X2=0.8910 $Y2=0.1530
r42 25 38 29.3819 $w=1.3e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.8125
+ $Y=0.1530 $X2=0.6865 $Y2=0.1530
r43 33 35 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.8910 $Y=0.1440
+ $X2=0.8910 $Y2=0.1530
r44 21 33 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1135 $X2=0.8910 $Y2=0.1440
r45 15 3 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.8910
+ $Y=0.1350 $X2=0.8910 $Y2=0.1350
r46 3 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8910 $Y=0.1350
+ $X2=0.8910 $Y2=0.1440
r47 8 17 1e-05
r48 7 16 1e-05
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%NET0120 VSS 13 24 26 8 1 2 9 11 10
c1 1 VSS 0.0056065f
c2 2 VSS 0.00858292f
c3 8 VSS 0.00327968f
c4 9 VSS 0.00235163f
c5 10 VSS 0.00214036f
c6 11 VSS 0.0211064f
r1 26 25 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r2 10 25 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5420 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r3 9 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4840 $Y2=0.2025
r4 24 9 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r5 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5130 $Y=0.2025
+ $X2=0.4900 $Y2=0.2340
r6 20 21 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4810
+ $Y=0.2340 $X2=0.4900 $Y2=0.2340
r7 19 20 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4690
+ $Y=0.2340 $X2=0.4810 $Y2=0.2340
r8 18 19 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4540
+ $Y=0.2340 $X2=0.4690 $Y2=0.2340
r9 17 18 17.7224 $w=1.3e-08 $l=7.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.4540 $Y2=0.2340
r10 16 17 19.5879 $w=1.3e-08 $l=8.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2940
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r11 15 16 5.59655 $w=1.3e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.2940 $Y2=0.2340
r12 11 15 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2580
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r13 8 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2160
+ $X2=0.2700 $Y2=0.2340
r14 1 8 23.8708 $w=2.02e-08 $l=4.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.2700 $Y=0.1755 $X2=0.2700 $Y2=0.2160
r15 13 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r16 8 12 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r17 2 10 1e-05
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%SI VSS 22 3 8 4 1 5 6 7
c1 1 VSS 0.00454521f
c2 3 VSS 0.0066463f
c3 4 VSS 0.00231197f
c4 5 VSS 0.00235282f
c5 6 VSS 0.00294562f
c6 7 VSS 0.00457396f
c7 8 VSS 0.00309483f
r1 6 21 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1980 $X2=0.5130 $Y2=0.1765
r2 23 24 5.65485 $w=1.3e-08 $l=2.43e-08 $layer=M2 $thickness=3.6e-08 $X=0.4887
+ $Y=0.1170 $X2=0.5130 $Y2=0.1170
r3 22 23 3.67274 $w=1.3e-08 $l=1.57e-08 $layer=M2 $thickness=3.6e-08 $X=0.4730
+ $Y=0.1170 $X2=0.4887 $Y2=0.1170
r4 22 8 0.757867 $w=1.3e-08 $l=3.3e-09 $layer=M2 $thickness=3.6e-08 $X=0.4730
+ $Y=0.1170 $X2=0.4697 $Y2=0.1170
r5 5 7 3.2503 $w=1.53684e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1540 $X2=0.5130 $Y2=0.1350
r6 5 21 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1540 $X2=0.5130 $Y2=0.1765
r7 20 24 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.5130 $Y=0.1170 $X2=0.5130
+ $Y2=0.1170
r8 7 18 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1350 $X2=0.4945 $Y2=0.1350
r9 7 20 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1170
r10 17 18 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4845
+ $Y=0.1350 $X2=0.4945 $Y2=0.1350
r11 16 17 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4750
+ $Y=0.1350 $X2=0.4845 $Y2=0.1350
r12 4 16 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4635
+ $Y=0.1350 $X2=0.4750 $Y2=0.1350
r13 14 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4790 $Y=0.1350
+ $X2=0.4750 $Y2=0.1350
r14 13 14 4.43042 $w=1.53e-08 $l=7.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.4715 $Y=0.1350 $X2=0.4790 $Y2=0.1350
r15 11 13 1.86855 $w=1.78125e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.4675 $Y=0.1350 $X2=0.4715 $Y2=0.1350
r16 1 11 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.4575
+ $Y=0.1350 $X2=0.4675 $Y2=0.1350
r17 3 1 2.53453 $w=1.32811e-07 $l=1.5e-09 $layer=LIG $thickness=5.23243e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4575 $Y2=0.1350
r18 3 13 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4715 $Y2=0.1350
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%PD5 VSS 7 12 4 1 5
c1 1 VSS 0.00743221f
c2 4 VSS 0.00187888f
c3 5 VSS 0.00236973f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9890 $Y=0.0405 $X2=0.9865 $Y2=0.0405
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9740 $Y=0.0405 $X2=0.9865 $Y2=0.0405
r3 9 5 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.9585
+ $Y=0.0405 $X2=0.9720 $Y2=0.0405
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.9435
+ $Y=0.0405 $X2=0.9585 $Y2=0.0405
r5 1 8 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.9180
+ $Y=0.0405 $X2=0.9435 $Y2=0.0405
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9035 $Y=0.0405 $X2=0.9160 $Y2=0.0405
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9010 $Y=0.0405 $X2=0.9035 $Y2=0.0405
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%PD3 VSS 2 4 1
c1 1 VSS 0.000910759f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.0405 $X2=0.7065 $Y2=0.0405
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.0405 $X2=0.6895 $Y2=0.0405
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6895 $Y=0.0405 $X2=0.7065 $Y2=0.0405
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%PD4 VSS 2 4 1
c1 1 VSS 0.00102278f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9890 $Y=0.2295 $X2=0.9765 $Y2=0.2295
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9550 $Y=0.2295 $X2=0.9595 $Y2=0.2295
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9595 $Y=0.2295 $X2=0.9765 $Y2=0.2295
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%noxref_26 VSS 1
c1 1 VSS 0.00432551f
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%PD2 VSS 7 12 4 5 1
c1 1 VSS 0.00742588f
c2 4 VSS 0.0018428f
c3 5 VSS 0.00234055f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7040 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r3 9 5 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.6765
+ $Y=0.2295 $X2=0.7020 $Y2=0.2295
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.6615
+ $Y=0.2295 $X2=0.6765 $Y2=0.2295
r5 1 8 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.6480
+ $Y=0.2295 $X2=0.6615 $Y2=0.2295
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.2295 $X2=0.6460 $Y2=0.2295
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.2295 $X2=0.6335 $Y2=0.2295
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%SS VSS 9 34 39 14 13 12 17 16 3 4 15 1 10 11
c1 1 VSS 0.00111365f
c2 3 VSS 0.00577733f
c3 4 VSS 0.00656554f
c4 9 VSS 0.0384079f
c5 10 VSS 0.00331732f
c6 11 VSS 0.00336502f
c7 12 VSS 0.00100028f
c8 13 VSS 0.00846082f
c9 14 VSS 0.00184799f
c10 15 VSS 0.00251824f
c11 16 VSS 0.00671548f
c12 17 VSS 0.0023068f
r1 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0655 $Y=0.2295 $X2=1.0780 $Y2=0.2295
r2 39 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0630 $Y=0.2295 $X2=1.0655 $Y2=0.2295
r3 4 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0800 $Y=0.2295
+ $X2=1.0800 $Y2=0.2340
r4 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.0800
+ $Y=0.2340 $X2=1.0935 $Y2=0.2340
r5 16 32 7.21452 $w=1.425e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.2340 $X2=1.1070 $Y2=0.1980
r6 16 37 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1070 $Y=0.2340 $X2=1.0935 $Y2=0.2340
r7 10 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.0655 $Y=0.0405 $X2=1.0780 $Y2=0.0405
r8 34 10 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.0630 $Y=0.0405 $X2=1.0655 $Y2=0.0405
r9 31 32 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.1440 $X2=1.1070 $Y2=0.1980
r10 14 30 8.95608 $w=1.36627e-08 $l=4.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1070 $Y=0.0810 $X2=1.1070 $Y2=0.0395
r11 14 31 14.691 $w=1.3e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.0810 $X2=1.1070 $Y2=0.1440
r12 3 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0800 $Y=0.0405
+ $X2=1.0800 $Y2=0.0360
r13 17 29 1.40651 $w=1.51875e-08 $l=1.45774e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1070 $Y=0.0305 $X2=1.0935 $Y2=0.0360
r14 17 30 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.0305 $X2=1.1070 $Y2=0.0395
r15 28 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.0800
+ $Y=0.0360 $X2=1.0935 $Y2=0.0360
r16 27 28 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.0685
+ $Y=0.0360 $X2=1.0800 $Y2=0.0360
r17 26 27 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.0640
+ $Y=0.0360 $X2=1.0685 $Y2=0.0360
r18 25 26 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.0360 $X2=1.0640 $Y2=0.0360
r19 13 15 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0260 $Y=0.0360 $X2=0.9990 $Y2=0.0360
r20 13 25 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.0360 $X2=1.0530 $Y2=0.0360
r21 12 22 8.04505 $w=1.3e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.9990
+ $Y=0.0705 $X2=0.9990 $Y2=0.1050
r22 12 15 6.39593 $w=1.55565e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9990 $Y=0.0705 $X2=0.9990 $Y2=0.0360
r23 1 19 2.36633 $w=2.3e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.9990
+ $Y=0.1055 $X2=0.9990 $Y2=0.1055
r24 1 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.9990 $Y=0.1055
+ $X2=0.9990 $Y2=0.1050
r25 9 19 0.314665 $w=2.27e-07 $l=2.95e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.9990 $Y=0.1350 $X2=0.9990 $Y2=0.1055
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%noxref_28 VSS 1
c1 1 VSS 0.00576953f
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%MS VSS 10 43 46 51 53 13 17 19 18 3 15 12 1 11 4
+ 14 16
c1 1 VSS 0.00318245f
c2 3 VSS 0.00574254f
c3 4 VSS 0.00955267f
c4 10 VSS 0.0376954f
c5 11 VSS 0.00302946f
c6 12 VSS 0.00287148f
c7 13 VSS 0.00239131f
c8 14 VSS 0.000902455f
c9 15 VSS 0.00367591f
c10 16 VSS 0.00188353f
c11 17 VSS 0.000914006f
c12 18 VSS 0.00131743f
c13 19 VSS 0.00120303f
c14 20 VSS 0.00289595f
r1 53 52 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8810 $Y=0.2295 $X2=0.8785 $Y2=0.2295
r2 13 52 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8660 $Y=0.2295 $X2=0.8785 $Y2=0.2295
r3 12 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.2295 $X2=0.8080 $Y2=0.2295
r4 51 12 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.2295 $X2=0.7955 $Y2=0.2295
r5 48 13 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8370 $Y=0.2295 $X2=0.8640 $Y2=0.2295
r6 4 48 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08 $X=0.8100
+ $Y=0.2295 $X2=0.8370 $Y2=0.2295
r7 4 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8100 $Y=0.2295
+ $X2=0.8125 $Y2=0.2340
r8 15 20 4.06404 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8125 $Y=0.2340 $X2=0.8370 $Y2=0.2340
r9 46 45 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8270 $Y=0.0405 $X2=0.8245 $Y2=0.0405
r10 44 45 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8200 $Y=0.0405 $X2=0.8245 $Y2=0.0405
r11 3 44 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8080 $Y=0.0405 $X2=0.8200 $Y2=0.0405
r12 11 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.0405 $X2=0.8080 $Y2=0.0405
r13 43 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.0405 $X2=0.7955 $Y2=0.0405
r14 20 39 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.2340 $X2=0.8370 $Y2=0.2160
r15 3 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8100 $Y=0.0405
+ $X2=0.8100 $Y2=0.0535
r16 38 39 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1870 $X2=0.8370 $Y2=0.2160
r17 37 38 4.89699 $w=1.3e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1660 $X2=0.8370 $Y2=0.1870
r18 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1525 $X2=0.8370 $Y2=0.1660
r19 35 36 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1310 $X2=0.8370 $Y2=0.1525
r20 34 35 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1115 $X2=0.8370 $Y2=0.1310
r21 17 31 1.15159 $w=1.75e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1000 $X2=0.8370 $Y2=0.0900
r22 17 34 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1000 $X2=0.8370 $Y2=0.1115
r23 16 32 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0625 $X2=0.8100 $Y2=0.0720
r24 16 33 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0625 $X2=0.8100 $Y2=0.0535
r25 30 31 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8235 $Y=0.0900 $X2=0.8370 $Y2=0.0900
r26 19 28 1.38478 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.0900 $X2=0.7990 $Y2=0.0900
r27 19 30 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.0900 $X2=0.8235 $Y2=0.0900
r28 19 32 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0900 $X2=0.8100 $Y2=0.0720
r29 27 28 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.7765
+ $Y=0.0900 $X2=0.7990 $Y2=0.0900
r30 14 27 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.7470
+ $Y=0.0900 $X2=0.7765 $Y2=0.0900
r31 14 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7470 $Y=0.0900
+ $X2=0.7500 $Y2=0.0900
r32 14 18 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7470
+ $Y=0.0900 $X2=0.7290 $Y2=0.0900
r33 25 26 5.02115 $w=1.53e-08 $l=8.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.7415 $Y=0.0900 $X2=0.7500 $Y2=0.0900
r34 23 25 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.7385 $Y=0.0900 $X2=0.7415 $Y2=0.0900
r35 1 23 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.7285
+ $Y=0.0900 $X2=0.7385 $Y2=0.0900
r36 1 22 2.48102 $w=2.2e-08 $l=5e-10 $layer=LIG $thickness=4.8e-08 $X=0.7285
+ $Y=0.0900 $X2=0.7290 $Y2=0.0900
r37 22 25 1.47681 $w=1.53e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7290 $Y=0.0900 $X2=0.7415 $Y2=0.0900
r38 10 22 0.314665 $w=2.27e-07 $l=4.5e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.7290 $Y=0.1350 $X2=0.7290 $Y2=0.0900
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%MH VSS 9 56 60 63 67 10 20 14 12 16 3 4 18 17 21
+ 1 19 15
c1 1 VSS 0.000205195f
c2 3 VSS 0.00474428f
c3 4 VSS 0.00497074f
c4 9 VSS 0.0362219f
c5 10 VSS 0.00228273f
c6 11 VSS 0.00010353f
c7 12 VSS 0.00212289f
c8 13 VSS 7.0661e-20
c9 14 VSS 0.00941548f
c10 15 VSS 0.00777258f
c11 16 VSS 0.00175484f
c12 17 VSS 0.000618516f
c13 18 VSS 0.00100604f
c14 19 VSS 0.00299202f
c15 20 VSS 5.91085e-20
c16 21 VSS 0.00269655f
r1 67 66 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.2295 $X2=0.6085 $Y2=0.2295
r2 65 66 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6040 $Y=0.2295 $X2=0.6085 $Y2=0.2295
r3 3 65 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5920 $Y=0.2295 $X2=0.6040 $Y2=0.2295
r4 13 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2295 $X2=0.5920 $Y2=0.2295
r5 61 62 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.1890 $X2=0.5840 $Y2=0.1890
r6 63 61 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.1890 $X2=0.5795 $Y2=0.1890
r7 12 62 0.185185 $w=5.4e-08 $l=1e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.1890 $X2=0.5840 $Y2=0.1890
r8 12 3 0.518519 $w=3.9e-08 $l=4.05494e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.1890 $X2=0.5920 $Y2=0.2295
r9 60 59 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r10 58 59 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6580 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r11 4 58 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6460 $Y=0.0405 $X2=0.6580 $Y2=0.0405
r12 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0405 $X2=0.6460 $Y2=0.0405
r13 10 4 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0810 $X2=0.6460 $Y2=0.0810
r14 56 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.0810 $X2=0.6335 $Y2=0.0810
r15 3 48 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2295
+ $X2=0.5900 $Y2=0.2340
r16 4 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.0405
+ $X2=0.6440 $Y2=0.0360
r17 45 46 1.63233 $w=1.3e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.5990
+ $Y=0.2340 $X2=0.6060 $Y2=0.2340
r18 45 48 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5990
+ $Y=0.2340 $X2=0.5900 $Y2=0.2340
r19 44 46 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.6105
+ $Y=0.2340 $X2=0.6060 $Y2=0.2340
r20 43 44 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6305
+ $Y=0.2340 $X2=0.6105 $Y2=0.2340
r21 14 21 4.53042 $w=1.46981e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6665 $Y=0.2340 $X2=0.6930 $Y2=0.2340
r22 14 43 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.6665
+ $Y=0.2340 $X2=0.6305 $Y2=0.2340
r23 15 40 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.6530
+ $Y=0.0360 $X2=0.6705 $Y2=0.0360
r24 15 42 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6530
+ $Y=0.0360 $X2=0.6440 $Y2=0.0360
r25 21 39 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.2340 $X2=0.6930 $Y2=0.2160
r26 19 34 2.43171 $w=1.804e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6930 $Y=0.0360 $X2=0.6930 $Y2=0.0535
r27 19 40 3.59766 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.0360 $X2=0.6705 $Y2=0.0360
r28 38 39 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1980 $X2=0.6930 $Y2=0.2160
r29 37 38 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1800 $X2=0.6930 $Y2=0.1980
r30 36 37 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1680 $X2=0.6930 $Y2=0.1800
r31 35 36 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1590 $X2=0.6930 $Y2=0.1680
r32 17 20 2.43413 $w=1.59032e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6930 $Y=0.1465 $X2=0.6930 $Y2=0.1310
r33 17 35 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1465 $X2=0.6930 $Y2=0.1590
r34 33 34 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.0625 $X2=0.6930 $Y2=0.0535
r35 32 33 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.0720 $X2=0.6930 $Y2=0.0625
r36 31 32 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.0900 $X2=0.6930 $Y2=0.0720
r37 30 31 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1025 $X2=0.6930 $Y2=0.0900
r38 16 20 2.78392 $w=1.56471e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6930 $Y=0.1140 $X2=0.6930 $Y2=0.1310
r39 16 30 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1140 $X2=0.6930 $Y2=0.1025
r40 20 28 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1310 $X2=0.7110 $Y2=0.1310
r41 27 28 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1310 $X2=0.7110 $Y2=0.1310
r42 18 26 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.1310 $X2=0.7830 $Y2=0.1310
r43 18 27 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.1310 $X2=0.7290 $Y2=0.1310
r44 1 23 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.7830
+ $Y=0.1310 $X2=0.7830 $Y2=0.1310
r45 1 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7830 $Y=0.1310
+ $X2=0.7830 $Y2=0.1310
r46 9 23 0.314665 $w=2.27e-07 $l=4e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.7830 $Y=0.1350 $X2=0.7830 $Y2=0.1310
r47 3 12 1e-05
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%noxref_27 VSS 1
c1 1 VSS 0.00430598f
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%noxref_29 VSS 1
c1 1 VSS 0.00584722f
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%noxref_30 VSS 1
c1 1 VSS 0.0126192f
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%NET0118 VSS 12 13 28 8 9 2 7 1
c1 1 VSS 0.00357752f
c2 2 VSS 0.00382155f
c3 7 VSS 0.00295314f
c4 8 VSS 0.00228056f
c5 9 VSS 0.00254762f
r1 28 27 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.0675 $X2=0.6085 $Y2=0.0675
r2 26 27 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6040 $Y=0.0675 $X2=0.6085 $Y2=0.0675
r3 8 26 0.123457 $w=8.1e-08 $l=1e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.0675 $X2=0.6040 $Y2=0.0675
r4 2 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0675
+ $X2=0.5900 $Y2=0.0720
r5 22 23 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.5805
+ $Y=0.0720 $X2=0.5900 $Y2=0.0720
r6 21 22 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0720 $X2=0.5805 $Y2=0.0720
r7 20 21 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.0720 $X2=0.5670 $Y2=0.0720
r8 19 20 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0720 $X2=0.5400 $Y2=0.0720
r9 18 19 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5020
+ $Y=0.0720 $X2=0.5130 $Y2=0.0720
r10 17 18 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4805
+ $Y=0.0720 $X2=0.5020 $Y2=0.0720
r11 16 17 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.4540
+ $Y=0.0720 $X2=0.4805 $Y2=0.0720
r12 15 16 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4440
+ $Y=0.0720 $X2=0.4540 $Y2=0.0720
r13 14 15 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0720 $X2=0.4440 $Y2=0.0720
r14 9 14 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4205
+ $Y=0.0720 $X2=0.4320 $Y2=0.0720
r15 1 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4320 $Y2=0.0720
r16 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r17 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r18 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0675 $X2=0.4320 $Y2=0.0675
r19 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4175 $Y2=0.0675
r20 2 8 1e-05
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%SE VSS 29 5 6 11 10 7 13 8 9 12 2 1
c1 1 VSS 0.00182947f
c2 2 VSS 0.00391123f
c3 5 VSS 0.0425749f
c4 6 VSS 0.0813612f
c5 7 VSS 0.00156595f
c6 8 VSS 0.000239343f
c7 9 VSS 0.00496752f
c8 10 VSS 0.00504547f
c9 11 VSS 0.000238173f
c10 12 VSS 0.00611557f
c11 13 VSS 0.0499567f
r1 1 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
r2 5 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r3 37 38 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2745
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r4 36 37 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2595
+ $Y=0.1350 $X2=0.2745 $Y2=0.1350
r5 35 36 0.699569 $w=1.3e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.1350 $X2=0.2595 $Y2=0.1350
r6 8 11 2.89809 $w=1.53077e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2445 $Y=0.1350 $X2=0.2250 $Y2=0.1350
r7 8 35 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2445
+ $Y=0.1350 $X2=0.2565 $Y2=0.1350
r8 11 33 3.59766 $w=1.692e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.1350 $X2=0.2250 $Y2=0.1125
r9 29 10 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.2250 $Y=0.0450 $X2=0.2250
+ $Y2=0.0360
r10 32 33 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0900 $X2=0.2250 $Y2=0.1125
r11 31 32 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0675 $X2=0.2250 $Y2=0.0900
r12 7 31 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0495 $X2=0.2250 $Y2=0.0675
r13 29 7 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.2250 $Y=0.0450 $X2=0.2250
+ $Y2=0.0495
r14 7 10 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.0495 $X2=0.2250 $Y2=0.0360
r15 29 30 7.92845 $w=1.3e-08 $l=3.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0450 $X2=0.2590 $Y2=0.0450
r16 27 30 12.0093 $w=1.3e-08 $l=5.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.3105
+ $Y=0.0450 $X2=0.2590 $Y2=0.0450
r17 26 27 103.886 $w=1.3e-08 $l=4.455e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.7560 $Y=0.0450 $X2=0.3105 $Y2=0.0450
r18 13 24 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=1.1905
+ $Y=0.0450 $X2=1.2150 $Y2=0.0450
r19 13 26 101.321 $w=1.3e-08 $l=4.345e-07 $layer=M2 $thickness=3.6e-08
+ $X=1.1905 $Y=0.0450 $X2=0.7560 $Y2=0.0450
r20 12 24 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=1.2150 $Y=0.0360 $X2=1.2150
+ $Y2=0.0450
r21 20 21 6.41272 $w=1.3e-08 $l=2.75e-08 $layer=M1 $thickness=3.6e-08 $X=1.2150
+ $Y=0.1085 $X2=1.2150 $Y2=0.1360
r22 19 20 8.51143 $w=1.3e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=1.2150
+ $Y=0.0720 $X2=1.2150 $Y2=0.1085
r23 9 19 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.2150
+ $Y=0.0495 $X2=1.2150 $Y2=0.0720
r24 9 12 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.2150 $Y=0.0495 $X2=1.2150 $Y2=0.0360
r25 9 24 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=1.2150 $Y=0.0495 $X2=1.2150
+ $Y2=0.0450
r26 6 2 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=1.2150
+ $Y=0.1350 $X2=1.2150 $Y2=0.1360
r27 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.2150 $Y=0.1360
+ $X2=1.2150 $Y2=0.1360
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%SH VSS 11 12 66 69 71 74 6 13 14 21 15 23 17 16 5
+ 25 20 2 22 1 18 19 24
c1 1 VSS 0.0006672f
c2 2 VSS 0.00367223f
c3 5 VSS 0.00496654f
c4 6 VSS 0.00511231f
c5 11 VSS 0.0378108f
c6 12 VSS 0.0800061f
c7 13 VSS 0.00364645f
c8 14 VSS 0.00383296f
c9 15 VSS 0.00797986f
c10 16 VSS 0.000578527f
c11 17 VSS 0.00136428f
c12 18 VSS 0.00118066f
c13 19 VSS 0.000154461f
c14 20 VSS 0.00335962f
c15 21 VSS 0.00653726f
c16 22 VSS 0.00216541f
c17 23 VSS 0.00010523f
c18 24 VSS 0.000358959f
c19 25 VSS 0.00991367f
r1 74 73 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8810 $Y=0.0405 $X2=0.8785 $Y2=0.0405
r2 5 73 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8660 $Y=0.0405 $X2=0.8785 $Y2=0.0405
r3 70 5 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8540 $Y=0.0405 $X2=0.8660 $Y2=0.0405
r4 13 70 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.0405 $X2=0.8540 $Y2=0.0405
r5 71 13 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.0405 $X2=0.8495 $Y2=0.0405
r6 69 68 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9350 $Y=0.2295 $X2=0.9325 $Y2=0.2295
r7 67 68 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9280 $Y=0.2295 $X2=0.9325 $Y2=0.2295
r8 6 67 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9160 $Y=0.2295 $X2=0.9280 $Y2=0.2295
r9 14 6 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9035 $Y=0.2295 $X2=0.9160 $Y2=0.2295
r10 66 14 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9010 $Y=0.2295 $X2=0.9035 $Y2=0.2295
r11 5 57 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.0405
+ $X2=0.8640 $Y2=0.0360
r12 6 52 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.9180 $Y=0.2295
+ $X2=0.9180 $Y2=0.2340
r13 2 49 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.2690 $Y=0.1360
+ $X2=1.2690 $Y2=0.1445
r14 12 2 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=1.2690
+ $Y=0.1350 $X2=1.2690 $Y2=0.1360
r15 57 58 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.0360 $X2=0.8775 $Y2=0.0360
r16 55 58 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.0360 $X2=0.8775 $Y2=0.0360
r17 54 55 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.9020
+ $Y=0.0360 $X2=0.8910 $Y2=0.0360
r18 15 22 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.9200
+ $Y=0.0360 $X2=0.9450 $Y2=0.0360
r19 15 54 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.9200
+ $Y=0.0360 $X2=0.9020 $Y2=0.0360
r20 52 53 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.2340 $X2=0.9315 $Y2=0.2340
r21 21 53 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.2340 $X2=0.9315 $Y2=0.2340
r22 20 49 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.2690
+ $Y=0.1085 $X2=1.2690 $Y2=0.1445
r23 22 43 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.0360 $X2=0.9450 $Y2=0.0630
r24 17 38 6.50021 $w=1.33448e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.1980 $X2=0.9450 $Y2=0.1690
r25 17 21 7.21452 $w=1.425e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.1980 $X2=0.9450 $Y2=0.2340
r26 47 49 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=1.2690 $Y=0.1530
+ $X2=1.2690 $Y2=0.1445
r27 46 47 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=1.2445
+ $Y=0.1530 $X2=1.2690 $Y2=0.1530
r28 45 46 9.91056 $w=1.3e-08 $l=4.25e-08 $layer=M2 $thickness=3.6e-08 $X=1.2020
+ $Y=0.1530 $X2=1.2445 $Y2=0.1530
r29 44 45 32.0636 $w=1.3e-08 $l=1.375e-07 $layer=M2 $thickness=3.6e-08
+ $X=1.0645 $Y=0.1530 $X2=1.2020 $Y2=0.1530
r30 25 44 27.8662 $w=1.3e-08 $l=1.195e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.9450 $Y=0.1530 $X2=1.0645 $Y2=0.1530
r31 25 39 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.9450 $Y=0.1530 $X2=0.9450
+ $Y2=0.1485
r32 42 43 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.0900 $X2=0.9450 $Y2=0.0630
r33 41 42 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1000 $X2=0.9450 $Y2=0.0900
r34 40 41 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1100 $X2=0.9450 $Y2=0.1000
r35 16 39 3.96423 $w=1.3e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1315 $X2=0.9450 $Y2=0.1485
r36 16 40 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1315 $X2=0.9450 $Y2=0.1100
r37 37 38 0.4592 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1645 $X2=0.9450 $Y2=0.1690
r38 23 37 0.714311 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1575 $X2=0.9450 $Y2=0.1645
r39 23 39 1.50855 $w=1.55e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1575 $X2=0.9450 $Y2=0.1485
r40 23 25 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.9450 $Y=0.1575 $X2=0.9450
+ $Y2=0.1530
r41 36 38 4.4015 $w=1.35e-08 $l=2.78927e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9720 $Y=0.1620 $X2=0.9450 $Y2=0.1690
r42 35 36 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9990
+ $Y=0.1620 $X2=0.9720 $Y2=0.1620
r43 18 24 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0260 $Y=0.1620 $X2=1.0530 $Y2=0.1620
r44 18 35 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.1620 $X2=0.9990 $Y2=0.1620
r45 24 33 0.915974 $w=2.10182e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0530 $Y=0.1620 $X2=1.0530 $Y2=0.1510
r46 32 33 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1400 $X2=1.0530 $Y2=0.1510
r47 19 32 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1250 $X2=1.0530 $Y2=0.1400
r48 1 29 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=1.0530
+ $Y=0.1400 $X2=1.0530 $Y2=0.1400
r49 1 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.0530 $Y=0.1400
+ $X2=1.0530 $Y2=0.1400
r50 11 29 0.314665 $w=2.27e-07 $l=5e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.0530 $Y=0.1350 $X2=1.0530 $Y2=0.1400
.ends

.subckt PM_SDFHx1_ASAP7_75t_R%CLKB VSS 14 15 16 17 85 87 19 20 18 26 7 6 23 24
+ 4 22 21 8 2 1 25
c1 1 VSS 0.000270688f
c2 2 VSS 6.58043e-20
c3 3 VSS 1e-36
c4 4 VSS 0.000292912f
c5 6 VSS 0.00736722f
c6 7 VSS 0.00737103f
c7 8 VSS 0.00382221f
c8 14 VSS 0.00584612f
c9 15 VSS 0.00509531f
c10 16 VSS 0.00438755f
c11 17 VSS 0.00518972f
c12 18 VSS 0.00773195f
c13 19 VSS 0.00766704f
c14 20 VSS 0.00331462f
c15 21 VSS 0.00131239f
c16 22 VSS 0.00134699f
c17 23 VSS 0.00581197f
c18 24 VSS 0.00579884f
c19 25 VSS 0.000596443f
c20 26 VSS 0.0248154f
r1 19 7 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1600 $Y2=0.2160
r2 87 19 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r3 18 6 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1600 $Y2=0.0540
r4 85 18 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r5 7 80 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r6 6 77 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r7 1 72 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1355
+ $X2=0.5670 $Y2=0.1350
r8 14 1 3.19489 $w=1.24e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1355
r9 80 81 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r10 24 68 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.1890 $Y2=0.2160
r11 24 81 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2340 $X2=0.1755 $Y2=0.2340
r12 77 78 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r13 23 65 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1890 $Y2=0.0630
r14 23 78 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1755 $Y2=0.0360
r15 25 69 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.1980 $X2=0.5670 $Y2=0.1845
r16 25 54 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.5670 $Y=0.1980 $X2=0.5670
+ $Y2=0.1890
r17 72 73 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1485
r18 70 73 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1620 $X2=0.5670 $Y2=0.1485
r19 21 69 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1755 $X2=0.5670 $Y2=0.1845
r20 21 70 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1755 $X2=0.5670 $Y2=0.1620
r21 67 68 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2025 $X2=0.1890 $Y2=0.2160
r22 66 67 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1935 $X2=0.1890 $Y2=0.2025
r23 64 65 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0900 $X2=0.1890 $Y2=0.0630
r24 63 64 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1100 $X2=0.1890 $Y2=0.0900
r25 62 63 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1325 $X2=0.1890 $Y2=0.1100
r26 61 62 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1540 $X2=0.1890 $Y2=0.1325
r27 60 61 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1655 $X2=0.1890 $Y2=0.1540
r28 58 59 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1735 $X2=0.1890 $Y2=0.1825
r29 58 60 1.86552 $w=1.3e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1735 $X2=0.1890 $Y2=0.1655
r30 20 59 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1870 $X2=0.1890 $Y2=0.1825
r31 20 66 1.51573 $w=1.3e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1870 $X2=0.1890 $Y2=0.1935
r32 55 56 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.6480
+ $Y=0.1890 $X2=0.7290 $Y2=0.1890
r33 54 55 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1890 $X2=0.6480 $Y2=0.1890
r34 54 69 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.5670 $Y=0.1890 $X2=0.5670
+ $Y2=0.1845
r35 53 54 44.0729 $w=1.3e-08 $l=1.89e-07 $layer=M2 $thickness=3.6e-08 $X=0.3780
+ $Y=0.1890 $X2=0.5670 $Y2=0.1890
r36 52 53 44.0729 $w=1.3e-08 $l=1.89e-07 $layer=M2 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1890 $X2=0.3780 $Y2=0.1890
r37 52 66 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1890 $Y=0.1890
+ $X2=0.1890 $Y2=0.1935
r38 26 52 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.1775
+ $Y=0.1890 $X2=0.1890 $Y2=0.1890
r39 4 49 2.78395 $w=2.4e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.9450
+ $Y=0.1780 $X2=0.9450 $Y2=0.1780
r40 17 4 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.9450 $Y=0.1350 $X2=0.9450 $Y2=0.1780
r41 2 42 2.78395 $w=2.4e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.6750
+ $Y=0.1780 $X2=0.6750 $Y2=0.1780
r42 15 2 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.6750 $Y=0.1350 $X2=0.6750 $Y2=0.1780
r43 50 56 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.7290 $Y=0.1845
+ $X2=0.7290 $Y2=0.1890
r44 22 50 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1680 $X2=0.7290 $Y2=0.1845
r45 48 49 6.83711 $w=2.22e-08 $l=1.5e-09 $layer=LISD $thickness=2.7e-08
+ $X=0.9435 $Y=0.1780 $X2=0.9450 $Y2=0.1780
r46 47 48 12.9145 $w=2.22e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9180 $Y=0.1780 $X2=0.9435 $Y2=0.1780
r47 46 47 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9045 $Y=0.1780 $X2=0.9180 $Y2=0.1780
r48 45 46 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8910 $Y=0.1780 $X2=0.9045 $Y2=0.1780
r49 44 45 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8775 $Y=0.1780 $X2=0.8910 $Y2=0.1780
r50 43 44 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8640 $Y=0.1780 $X2=0.8775 $Y2=0.1780
r51 41 42 12.9145 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6885 $Y=0.1780 $X2=0.6750 $Y2=0.1780
r52 40 41 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7155 $Y=0.1780 $X2=0.6885 $Y2=0.1780
r53 38 39 6.07743 $w=2.22e-08 $l=1.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7290 $Y=0.1780 $X2=0.7410 $Y2=0.1780
r54 38 50 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7290 $Y=0.1780
+ $X2=0.7290 $Y2=0.1845
r55 37 38 5.31775 $w=2.22e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7185 $Y=0.1780 $X2=0.7290 $Y2=0.1780
r56 37 40 1.51936 $w=2.22e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.7185
+ $Y=0.1780 $X2=0.7155 $Y2=0.1780
r57 36 39 4.55807 $w=2.22e-08 $l=9e-09 $layer=LISD $thickness=2.7e-08 $X=0.7500
+ $Y=0.1780 $X2=0.7410 $Y2=0.1780
r58 35 36 6.07743 $w=2.22e-08 $l=1.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7620 $Y=0.1780 $X2=0.7500 $Y2=0.1780
r59 34 35 4.05162 $w=2.22e-08 $l=8e-09 $layer=LISD $thickness=2.7e-08 $X=0.7700
+ $Y=0.1780 $X2=0.7620 $Y2=0.1780
r60 33 34 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7835 $Y=0.1780 $X2=0.7700 $Y2=0.1780
r61 32 33 6.58388 $w=2.22e-08 $l=1.3e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7965 $Y=0.1780 $X2=0.7835 $Y2=0.1780
r62 31 32 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8100 $Y=0.1780 $X2=0.7965 $Y2=0.1780
r63 8 31 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8370 $Y=0.1780 $X2=0.8100 $Y2=0.1780
r64 8 43 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8370 $Y=0.1780 $X2=0.8640 $Y2=0.1780
r65 3 30 2.78395 $w=2.4e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.8370
+ $Y=0.1780 $X2=0.8370 $Y2=0.1780
r66 3 8 10.3807 $w=2.30357e-08 $l=0 $layer=LISD $thickness=3.675e-08 $X=0.8370
+ $Y=0.1780 $X2=0.8370 $Y2=0.1780
r67 16 30 0.314665 $w=2.27e-07 $l=4.3e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.8370 $Y=0.1350 $X2=0.8370 $Y2=0.1780
.ends


*
.SUBCKT SDFHx1_ASAP7_75t_R VSS VDD CLK SE D SI QN
*
* VSS VSS
* VDD VDD
* CLK CLK
* SE SE
* D D
* SI SI
* QN QN
*
*

MM20 N_MM20_d N_MM20_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM23 N_MM23_d N_MM22_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM0 N_MM0_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM28 N_MM28_d N_MM2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM29 N_MM29_d N_MM26_g N_MM29_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM27_g N_MM5_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM10_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM6 N_MM6_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM12 N_MM12_d N_MM12_g N_MM12_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM17 N_MM17_d N_MM17_g N_MM17_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM16 N_MM16_d N_MM16_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM14 N_MM14_d N_MM14_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM30 N_MM30_d N_MM30_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM24 N_MM24_d N_MM24_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM21 N_MM21_d N_MM20_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM22 N_MM22_d N_MM22_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g N_MM3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM26 N_MM26_d N_MM26_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM27 N_MM27_d N_MM27_g N_MM27_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM13 N_MM13_d N_MM17_g N_MM13_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM18 N_MM18_d N_MM18_g N_MM18_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM19 N_MM19_d N_MM16_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM15 N_MM15_d N_MM14_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM31 N_MM31_d N_MM30_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM25 N_MM25_d N_MM24_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "SDFHx1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "SDFHx1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_SDFHx1_ASAP7_75t_R%NET0166 VSS N_MM28_d N_MM29_s N_NET0166_1
+ PM_SDFHx1_ASAP7_75t_R%NET0166
cc_1 N_NET0166_1 N_MM2_g 0.0173497f
cc_2 N_NET0166_1 N_MM26_g 0.0172412f
x_PM_SDFHx1_ASAP7_75t_R%noxref_31 VSS N_noxref_31_1
+ PM_SDFHx1_ASAP7_75t_R%noxref_31
cc_3 N_noxref_31_1 N_SEN_3 0.00118547f
cc_4 N_noxref_31_1 N_SS_10 0.0170009f
cc_5 N_noxref_31_1 N_MM14_g 0.00574621f
x_PM_SDFHx1_ASAP7_75t_R%noxref_32 VSS N_noxref_32_1
+ PM_SDFHx1_ASAP7_75t_R%noxref_32
cc_6 N_noxref_32_1 N_SEN_11 0.000619391f
cc_7 N_noxref_32_1 N_SS_11 0.0170395f
cc_8 N_noxref_32_1 N_MM14_g 0.00582034f
cc_9 N_noxref_32_1 N_noxref_31_1 0.00153605f
x_PM_SDFHx1_ASAP7_75t_R%noxref_33 VSS N_noxref_33_1
+ PM_SDFHx1_ASAP7_75t_R%noxref_33
cc_10 N_noxref_33_1 N_MM30_g 0.00558924f
cc_11 N_noxref_33_1 N_SEN_3 0.00143457f
cc_12 N_noxref_33_1 N_SEN_10 0.0170343f
cc_13 N_noxref_33_1 N_SS_10 0.000444701f
cc_14 N_noxref_33_1 N_noxref_31_1 0.00768437f
cc_15 N_noxref_33_1 N_noxref_32_1 0.000508626f
x_PM_SDFHx1_ASAP7_75t_R%noxref_34 VSS N_noxref_34_1
+ PM_SDFHx1_ASAP7_75t_R%noxref_34
cc_16 N_noxref_34_1 N_SE_2 0.000170279f
cc_17 N_noxref_34_1 N_MM30_g 0.00552392f
cc_18 N_noxref_34_1 N_SEN_13 0.000207857f
cc_19 N_noxref_34_1 N_SEN_4 0.000300559f
cc_20 N_noxref_34_1 N_SEN_11 0.0164753f
cc_21 N_noxref_34_1 N_SS_11 0.000611892f
cc_22 N_noxref_34_1 N_noxref_31_1 0.000510561f
cc_23 N_noxref_34_1 N_noxref_32_1 0.0078672f
cc_24 N_noxref_34_1 N_noxref_33_1 0.00152564f
x_PM_SDFHx1_ASAP7_75t_R%NET0167 VSS N_MM0_d N_MM5_s N_NET0167_7 N_NET0167_9
+ N_NET0167_1 N_NET0167_11 N_NET0167_12 N_NET0167_10 N_NET0167_8 N_NET0167_2
+ PM_SDFHx1_ASAP7_75t_R%NET0167
cc_25 N_NET0167_7 N_SE_1 0.00126965f
cc_26 N_NET0167_9 N_SE_10 0.000751402f
cc_27 N_NET0167_1 N_SE_8 0.000835429f
cc_28 N_NET0167_11 N_SE_7 0.00128783f
cc_29 N_NET0167_12 N_SE_10 0.00131201f
cc_30 N_NET0167_1 N_MM3_g 0.00158822f
cc_31 N_NET0167_11 N_SE_8 0.00339766f
cc_32 N_NET0167_10 N_SE_13 0.00420573f
cc_33 N_NET0167_7 N_MM3_g 0.0341503f
cc_34 N_NET0167_10 N_SEN_12 0.000311072f
cc_35 N_NET0167_10 N_SEN_16 0.000322875f
cc_36 N_NET0167_11 N_SEN_12 0.00107706f
cc_37 N_NET0167_10 N_SEN_14 0.00522531f
cc_38 N_NET0167_8 N_SI_1 0.00130085f
cc_39 N_NET0167_2 N_MM27_g 0.0015411f
cc_40 N_NET0167_8 N_MM27_g 0.0348642f
x_PM_SDFHx1_ASAP7_75t_R%noxref_35 VSS N_noxref_35_1
+ PM_SDFHx1_ASAP7_75t_R%noxref_35
cc_41 N_noxref_35_1 N_MM24_g 0.00147581f
cc_42 N_noxref_35_1 N_QN_7 0.038496f
x_PM_SDFHx1_ASAP7_75t_R%noxref_36 VSS N_noxref_36_1
+ PM_SDFHx1_ASAP7_75t_R%noxref_36
cc_43 N_noxref_36_1 N_MM24_g 0.00147666f
cc_44 N_noxref_36_1 N_QN_8 0.0384392f
cc_45 N_noxref_36_1 N_noxref_35_1 0.00176716f
x_PM_SDFHx1_ASAP7_75t_R%QN VSS QN N_MM24_d N_MM25_d N_QN_10 N_QN_7 N_QN_11
+ N_QN_2 N_QN_1 N_QN_8 N_QN_9 PM_SDFHx1_ASAP7_75t_R%QN
cc_46 N_QN_10 N_SE_9 0.000786105f
cc_47 N_QN_10 N_SE_13 0.00024607f
cc_48 N_QN_10 N_SE_12 0.00164048f
cc_49 N_QN_7 N_SH_20 0.00124847f
cc_50 N_QN_11 N_SH_25 0.000705726f
cc_51 N_QN_2 N_SH_2 0.000753967f
cc_52 N_QN_1 N_MM24_g 0.00119711f
cc_53 N_QN_2 N_MM24_g 0.00137744f
cc_54 N_QN_8 N_SH_2 0.00173173f
cc_55 N_QN_8 N_MM24_g 0.0150939f
cc_56 N_QN_9 N_SH_20 0.00674891f
cc_57 N_QN_7 N_MM24_g 0.0545134f
x_PM_SDFHx1_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_SDFHx1_ASAP7_75t_R%noxref_25
cc_58 N_noxref_25_1 N_MM20_g 0.00368844f
cc_59 N_noxref_25_1 N_CLKN_23 5.55503e-20
cc_60 N_noxref_25_1 N_CLKN_18 0.000383509f
cc_61 N_noxref_25_1 N_CLKN_8 0.000504425f
cc_62 N_noxref_25_1 N_CLKN_17 0.0275425f
cc_63 N_noxref_25_1 N_noxref_24_1 0.00204604f
x_PM_SDFHx1_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_SDFHx1_ASAP7_75t_R%noxref_24
cc_64 N_noxref_24_1 N_MM20_g 0.00366986f
cc_65 N_noxref_24_1 N_CLKN_22 5.93557e-20
cc_66 N_noxref_24_1 N_CLKN_18 0.000385062f
cc_67 N_noxref_24_1 N_CLKN_7 0.000429768f
cc_68 N_noxref_24_1 N_CLKN_16 0.0275836f
x_PM_SDFHx1_ASAP7_75t_R%D VSS D N_MM26_g N_D_5 N_D_4 N_D_1
+ PM_SDFHx1_ASAP7_75t_R%D
cc_69 N_D_5 N_CLKN_25 0.0139564f
cc_70 N_D_5 N_SE_8 0.000306664f
cc_71 N_D_5 N_SE_13 0.00240076f
cc_72 N_D_5 N_SEN_14 0.000401754f
cc_73 N_D_5 N_SEN_12 0.000468639f
cc_74 N_D_4 N_SEN_16 0.000640871f
cc_75 N_D_1 N_SEN_1 0.00211518f
cc_76 N_D_4 N_SEN_12 0.00286507f
cc_77 N_MM26_g N_MM2_g 0.00498026f
cc_78 N_D_5 N_SEN_16 0.00891151f
x_PM_SDFHx1_ASAP7_75t_R%SEN VSS N_MM2_g N_MM30_d N_MM31_d N_SEN_16 N_SEN_12
+ N_SEN_14 N_SEN_4 N_SEN_10 N_SEN_11 N_SEN_13 N_SEN_3 N_SEN_1 N_SEN_15
+ PM_SDFHx1_ASAP7_75t_R%SEN
cc_79 N_SEN_16 N_CLKN_21 0.00307496f
cc_80 N_SEN_16 N_CLKN_20 0.000328408f
cc_81 N_SEN_12 N_CLKN_25 0.00123727f
cc_82 N_SEN_16 N_CLKN_25 0.00662623f
cc_83 N_SEN_14 N_SE_13 0.000209557f
cc_84 N_SEN_4 N_SE_9 0.000213964f
cc_85 N_SEN_10 N_MM30_g 0.0232234f
cc_86 N_SEN_11 N_MM30_g 0.00679662f
cc_87 N_SEN_13 N_SE_9 0.00795256f
cc_88 N_SEN_3 N_SE_9 0.000259952f
cc_89 N_SEN_1 N_SE_8 0.0002982f
cc_90 N_SEN_13 N_SE_12 0.000329558f
cc_91 N_SEN_4 N_MM30_g 0.000349196f
cc_92 N_SEN_13 N_SE_2 0.000398285f
cc_93 N_SEN_3 N_SE_2 0.000413442f
cc_94 N_SEN_15 N_SE_9 0.000417695f
cc_95 N_SEN_1 N_SE_1 0.00129004f
cc_96 N_SEN_12 N_SE_13 0.000453145f
cc_97 N_SEN_13 N_SE_13 0.000514998f
cc_98 N_SEN_3 N_MM30_g 0.00098246f
cc_99 N_SEN_12 N_SE_8 0.00164495f
cc_100 N_MM2_g N_MM3_g 0.00330889f
cc_101 N_SEN_16 N_SE_13 0.0621894f
x_PM_SDFHx1_ASAP7_75t_R%CLK VSS CLK N_MM20_g N_CLK_6 N_CLK_8 N_CLK_1 N_CLK_5
+ N_CLK_4 N_CLK_7 PM_SDFHx1_ASAP7_75t_R%CLK
x_PM_SDFHx1_ASAP7_75t_R%NET0141 VSS N_MM3_s N_MM2_d N_MM26_d N_MM27_s
+ N_NET0141_7 N_NET0141_9 N_NET0141_1 N_NET0141_8 N_NET0141_2
+ PM_SDFHx1_ASAP7_75t_R%NET0141
cc_102 N_NET0141_7 N_SE_1 0.00103169f
cc_103 N_NET0141_9 N_SE_8 0.000641102f
cc_104 N_NET0141_1 N_MM3_g 0.000835657f
cc_105 N_NET0141_7 N_MM3_g 0.0329441f
cc_106 N_NET0141_7 N_SEN_1 0.000918818f
cc_107 N_NET0141_1 N_MM2_g 0.000852341f
cc_108 N_NET0141_9 N_SEN_12 0.00219558f
cc_109 N_NET0141_7 N_MM2_g 0.0329903f
cc_110 N_NET0141_8 N_D_1 0.000589038f
cc_111 N_NET0141_2 N_MM26_g 0.000900338f
cc_112 N_NET0141_9 N_D_4 0.00231406f
cc_113 N_NET0141_8 N_MM26_g 0.033409f
cc_114 N_NET0141_9 N_SI_4 0.000702864f
cc_115 N_NET0141_8 N_SI_1 0.000778696f
cc_116 N_NET0141_2 N_MM27_g 0.00083423f
cc_117 N_NET0141_8 N_MM27_g 0.0335665f
cc_118 N_NET0141_9 N_CLKB_26 0.00301772f
cc_119 N_NET0141_2 N_NET0120_11 0.000548369f
cc_120 N_NET0141_7 N_NET0120_8 0.00110519f
cc_121 N_NET0141_8 N_NET0120_9 0.000554907f
cc_122 N_NET0141_1 N_NET0120_11 0.000597641f
cc_123 N_NET0141_8 N_NET0120_2 0.00130017f
cc_124 N_NET0141_2 N_NET0120_2 0.00160616f
cc_125 N_NET0141_1 N_NET0120_1 0.00303079f
cc_126 N_NET0141_9 N_NET0120_11 0.0130912f
x_PM_SDFHx1_ASAP7_75t_R%CLKN VSS N_MM22_g N_MM10_g N_MM17_g N_MM20_d N_MM21_d
+ N_CLKN_8 N_CLKN_18 N_CLKN_7 N_CLKN_17 N_CLKN_16 N_CLKN_19 N_CLKN_1 N_CLKN_23
+ N_CLKN_25 N_CLKN_22 N_CLKN_21 N_CLKN_20 N_CLKN_3 N_CLKN_2 N_CLKN_24
+ PM_SDFHx1_ASAP7_75t_R%CLKN
cc_127 N_CLKN_8 N_MM20_g 0.00108708f
cc_128 N_CLKN_18 N_MM20_g 0.000251584f
cc_129 N_CLKN_7 N_MM20_g 0.00110453f
cc_130 N_CLKN_17 N_MM20_g 0.0112174f
cc_131 N_CLKN_16 N_MM20_g 0.0112195f
cc_132 N_CLKN_19 N_MM20_g 0.00034984f
cc_133 N_CLKN_1 N_CLK_6 0.000709538f
cc_134 N_CLKN_23 N_CLK_8 0.000822621f
cc_135 N_CLKN_19 N_CLK_8 0.000893482f
cc_136 N_CLKN_1 N_CLK_1 0.0034236f
cc_137 N_CLKN_18 N_CLK_6 0.000951613f
cc_138 N_CLKN_19 N_CLK_6 0.00105675f
cc_139 N_CLKN_25 N_CLK_8 0.00154373f
cc_140 N_CLKN_22 N_CLK_5 0.00172794f
cc_141 N_CLKN_19 N_CLK_4 0.00174141f
cc_142 N_CLKN_23 N_CLK_7 0.0019618f
cc_143 N_CLKN_18 N_CLK_4 0.00658767f
cc_144 N_MM22_g N_MM20_g 0.035014f
x_PM_SDFHx1_ASAP7_75t_R%NET0120 VSS N_MM3_d N_MM27_d N_MM1_s N_NET0120_8
+ N_NET0120_1 N_NET0120_2 N_NET0120_9 N_NET0120_11 N_NET0120_10
+ PM_SDFHx1_ASAP7_75t_R%NET0120
cc_145 N_NET0120_8 N_SE_11 0.000124442f
cc_146 N_NET0120_8 N_SE_8 0.000691325f
cc_147 N_NET0120_8 N_SE_1 0.00106117f
cc_148 N_NET0120_1 N_MM3_g 0.00131448f
cc_149 N_NET0120_8 N_MM3_g 0.0339702f
cc_150 N_NET0120_2 N_SI_5 0.000637517f
cc_151 N_NET0120_9 N_SI_1 0.00143551f
cc_152 N_NET0120_2 N_SI_6 0.00293538f
cc_153 N_NET0120_11 N_SI_6 0.00311408f
cc_154 N_NET0120_9 N_MM27_g 0.0349925f
cc_155 N_NET0120_10 N_CLKB_20 4.84051e-20
cc_156 N_NET0120_10 N_CLKB_24 0.000288049f
cc_157 N_NET0120_10 N_CLKB_7 0.000136682f
cc_158 N_NET0120_10 N_CLKB_19 0.000143172f
cc_159 N_NET0120_10 N_CLKB_1 0.00101238f
cc_160 N_NET0120_10 N_CLKB_25 0.000340224f
cc_161 N_NET0120_10 N_CLKB_21 0.00035735f
cc_162 N_NET0120_1 N_CLKB_20 0.000942542f
cc_163 N_NET0120_2 N_MM1_g 0.00158906f
cc_164 N_NET0120_11 N_CLKB_26 0.00353064f
cc_165 N_NET0120_10 N_MM1_g 0.0338896f
cc_166 N_NET0120_2 N_MH_3 0.00118806f
cc_167 N_NET0120_2 N_MH_12 0.00291444f
x_PM_SDFHx1_ASAP7_75t_R%SI VSS SI N_MM27_g N_SI_8 N_SI_4 N_SI_1 N_SI_5 N_SI_6
+ N_SI_7 PM_SDFHx1_ASAP7_75t_R%SI
cc_168 N_SI_8 N_CLKN_20 0.000103317f
cc_169 N_SI_4 N_CLKN_25 0.000849835f
cc_170 N_SI_8 N_CLKN_25 0.0114174f
cc_171 N_SI_8 N_SEN_16 0.0104368f
cc_172 N_SI_8 N_MM26_g 0.000739684f
cc_173 N_SI_1 N_D_1 0.000866384f
cc_174 N_SI_4 N_D_4 0.000945027f
cc_175 N_MM27_g N_MM26_g 0.00377702f
x_PM_SDFHx1_ASAP7_75t_R%PD5 VSS N_MM17_s N_MM16_d N_PD5_4 N_PD5_1 N_PD5_5
+ PM_SDFHx1_ASAP7_75t_R%PD5
cc_176 N_PD5_4 N_CLKN_3 9.95216e-20
cc_177 N_PD5_4 N_MM17_g 0.0151527f
cc_178 N_PD5_1 N_MM18_g 0.000757468f
cc_179 N_PD5_5 N_MM18_g 0.00693206f
cc_180 N_PD5_4 N_MM18_g 0.0239763f
cc_181 N_PD5_1 N_MM16_g 0.000891908f
cc_182 N_PD5_5 N_MM16_g 0.0155917f
cc_183 N_PD5_1 N_SH_13 0.000514787f
cc_184 N_PD5_1 N_SH_15 0.000490359f
cc_185 N_PD5_1 N_SH_16 0.000570793f
cc_186 N_PD5_4 N_SH_5 0.000657964f
cc_187 N_PD5_1 N_SH_22 0.00237801f
x_PM_SDFHx1_ASAP7_75t_R%PD3 VSS N_MM9_s N_MM8_d N_PD3_1
+ PM_SDFHx1_ASAP7_75t_R%PD3
cc_188 N_PD3_1 N_MM9_g 0.00777458f
cc_189 N_PD3_1 N_MM11_g 0.00783316f
x_PM_SDFHx1_ASAP7_75t_R%PD4 VSS N_MM18_s N_MM19_d N_PD4_1
+ PM_SDFHx1_ASAP7_75t_R%PD4
cc_190 N_PD4_1 N_MM18_g 0.00783925f
cc_191 N_PD4_1 N_MM16_g 0.00773636f
x_PM_SDFHx1_ASAP7_75t_R%noxref_26 VSS N_noxref_26_1
+ PM_SDFHx1_ASAP7_75t_R%noxref_26
cc_192 N_noxref_26_1 N_MM22_g 0.00351507f
cc_193 N_noxref_26_1 N_CLKB_20 0.000145915f
cc_194 N_noxref_26_1 N_CLKB_6 0.000432466f
cc_195 N_noxref_26_1 N_CLKB_18 0.0270445f
cc_196 N_noxref_26_1 N_NET0167_7 0.00055795f
x_PM_SDFHx1_ASAP7_75t_R%PD2 VSS N_MM10_s N_MM11_d N_PD2_4 N_PD2_5 N_PD2_1
+ PM_SDFHx1_ASAP7_75t_R%PD2
cc_197 N_PD2_4 N_MM10_g 0.0150121f
cc_198 N_PD2_4 N_CLKB_8 0.000122246f
cc_199 N_PD2_4 N_CLKB_2 0.000277556f
cc_200 N_PD2_5 N_CLKB_8 0.00167232f
cc_201 N_PD2_1 N_MM9_g 0.00209541f
cc_202 N_PD2_5 N_MM9_g 0.0073462f
cc_203 N_PD2_4 N_MM9_g 0.0238309f
cc_204 N_PD2_5 N_MM11_g 0.0148527f
cc_205 N_PD2_4 N_MH_14 0.000321585f
cc_206 N_PD2_1 N_MH_17 0.000354751f
cc_207 N_PD2_4 N_MH_3 0.000612778f
cc_208 N_PD2_1 N_MH_14 0.0031281f
x_PM_SDFHx1_ASAP7_75t_R%SS VSS N_MM16_g N_MM14_d N_MM15_d N_SS_14 N_SS_13
+ N_SS_12 N_SS_17 N_SS_16 N_SS_3 N_SS_4 N_SS_15 N_SS_1 N_SS_10 N_SS_11
+ PM_SDFHx1_ASAP7_75t_R%SS
cc_209 N_SS_14 N_SE_13 0.000526247f
cc_210 N_SS_13 N_SE_13 0.000906364f
cc_211 N_SS_12 N_SE_13 0.00292927f
cc_212 N_SS_14 N_SEN_3 0.00127833f
cc_213 N_SS_14 N_SEN_4 0.000106965f
cc_214 N_SS_14 N_SEN_15 0.000108856f
cc_215 N_SS_13 N_SEN_16 0.00035578f
cc_216 N_SS_17 N_SEN_13 0.000424246f
cc_217 N_SS_16 N_SEN_15 0.000788213f
cc_218 N_SS_12 N_SEN_16 0.00260718f
cc_219 N_SS_14 N_SEN_13 0.00825663f
cc_220 N_MM16_g N_CLKB_8 0.000681186f
cc_221 N_MM16_g N_CLKB_4 0.000426619f
cc_222 N_MM16_g N_MM18_g 0.0133451f
x_PM_SDFHx1_ASAP7_75t_R%noxref_28 VSS N_noxref_28_1
+ PM_SDFHx1_ASAP7_75t_R%noxref_28
cc_223 N_noxref_28_1 N_MM3_g 0.00164816f
cc_224 N_noxref_28_1 N_CLKB_6 9.95924e-20
cc_225 N_noxref_28_1 N_CLKB_18 0.000515035f
cc_226 N_noxref_28_1 N_NET0167_7 0.0359949f
cc_227 N_noxref_28_1 N_noxref_26_1 0.00769512f
cc_228 N_noxref_28_1 N_noxref_27_1 0.00046973f
x_PM_SDFHx1_ASAP7_75t_R%MS VSS N_MM11_g N_MM6_d N_MM12_d N_MM7_d N_MM13_d
+ N_MS_13 N_MS_17 N_MS_19 N_MS_18 N_MS_3 N_MS_15 N_MS_12 N_MS_1 N_MS_11 N_MS_4
+ N_MS_14 N_MS_16 PM_SDFHx1_ASAP7_75t_R%MS
cc_229 N_MS_13 N_CLKN_21 0.0002466f
cc_230 N_MS_13 N_MM10_g 0.000137901f
cc_231 N_MS_13 N_CLKN_25 0.000344534f
cc_232 N_MS_13 N_CLKN_3 0.000222252f
cc_233 N_MS_17 N_CLKN_21 0.00432973f
cc_234 N_MS_17 N_CLKN_3 0.000289706f
cc_235 N_MS_19 N_CLKN_21 0.000412165f
cc_236 N_MS_18 N_CLKN_25 0.00159353f
cc_237 N_MS_13 N_MM17_g 0.0155043f
cc_238 N_MS_18 N_SEN_16 0.000904569f
cc_239 N_MS_19 N_SEN_16 0.00298001f
cc_240 N_MS_3 N_CLKB_22 0.000141461f
cc_241 N_MS_3 N_CLKB_8 0.000630961f
cc_242 N_MS_3 N_CLKB_2 9.2565e-20
cc_243 N_MS_3 N_CLKB_26 0.000143017f
cc_244 N_MS_15 N_CLKB_22 0.000275964f
cc_245 N_MS_13 N_MM12_g 0.00786932f
cc_246 N_MS_12 N_MM12_g 0.00781542f
cc_247 N_MS_15 N_CLKB_8 0.000372105f
cc_248 N_MS_1 N_MM9_g 0.000704085f
cc_249 N_MS_17 N_CLKB_8 0.00159528f
cc_250 N_MS_11 N_MM12_g 0.00650899f
cc_251 N_MS_4 N_MM12_g 0.002572f
cc_252 N_MS_4 N_CLKB_8 0.00638415f
cc_253 N_MM11_g N_MM9_g 0.014171f
cc_254 N_MS_3 N_MM12_g 0.0259928f
x_PM_SDFHx1_ASAP7_75t_R%MH VSS N_MM7_g N_MM4_d N_MM9_d N_MM1_d N_MM10_d N_MH_10
+ N_MH_20 N_MH_14 N_MH_12 N_MH_16 N_MH_3 N_MH_4 N_MH_18 N_MH_17 N_MH_21 N_MH_1
+ N_MH_19 N_MH_15 PM_SDFHx1_ASAP7_75t_R%MH
cc_255 N_MH_10 N_CLKN_3 0.00010891f
cc_256 N_MH_10 N_CLKN_20 0.000254717f
cc_257 N_MH_10 N_MM17_g 0.000137198f
cc_258 N_MH_10 N_CLKN_24 0.000294355f
cc_259 N_MH_20 N_CLKN_24 0.00031833f
cc_260 N_MH_14 N_CLKN_24 0.000444103f
cc_261 N_MH_12 N_MM10_g 0.0163939f
cc_262 N_MH_16 N_CLKN_20 0.000524098f
cc_263 N_MH_3 N_CLKN_2 0.000605753f
cc_264 N_MH_4 N_CLKN_20 0.000780464f
cc_265 N_MH_18 N_CLKN_25 0.000956505f
cc_266 N_MH_4 N_MM10_g 0.00111259f
cc_267 N_MH_3 N_MM10_g 0.00122592f
cc_268 N_MH_10 N_CLKN_2 0.00161087f
cc_269 N_MH_17 N_CLKN_25 0.00164425f
cc_270 N_MH_17 N_CLKN_24 0.0020624f
cc_271 N_MH_10 N_MM10_g 0.0527673f
cc_272 N_MH_10 N_CLKB_21 0.00012253f
cc_273 N_MH_10 N_CLKB_22 0.000340744f
cc_274 N_MH_10 N_MM1_g 0.000428971f
cc_275 N_MH_10 N_CLKB_1 0.000203325f
cc_276 N_MH_3 N_CLKB_21 0.000351862f
cc_277 N_MH_3 N_CLKB_25 0.000359961f
cc_278 N_MH_21 N_CLKB_22 0.000404645f
cc_279 N_MH_17 N_CLKB_22 0.00611995f
cc_280 N_MH_17 N_CLKB_2 0.000498197f
cc_281 N_MH_1 N_CLKB_8 0.00211257f
cc_282 N_MH_4 N_MM9_g 0.00063453f
cc_283 N_MH_12 N_CLKB_1 0.000668692f
cc_284 N_MH_17 N_CLKB_8 0.000742732f
cc_285 N_MH_14 N_CLKB_26 0.00140508f
cc_286 N_MH_18 N_CLKB_22 0.00148898f
cc_287 N_MH_3 N_MM1_g 0.00156549f
cc_288 N_MH_14 N_CLKB_25 0.00378042f
cc_289 N_MM7_g N_CLKB_8 0.00510582f
cc_290 N_MH_12 N_MM1_g 0.0330337f
cc_291 N_MM7_g N_MM12_g 0.0127578f
cc_292 N_MH_10 N_MM9_g 0.0362197f
cc_293 N_MH_19 N_MS_18 0.000267655f
cc_294 N_MH_4 N_MS_1 0.000360935f
cc_295 N_MH_18 N_MS_19 0.000419775f
cc_296 N_MH_18 N_MS_1 0.000676175f
cc_297 N_MH_1 N_MS_14 0.000871573f
cc_298 N_MM7_g N_MS_3 0.000940779f
cc_299 N_MH_18 N_MS_17 0.000984691f
cc_300 N_MH_1 N_MS_1 0.00130665f
cc_301 N_MM7_g N_MS_12 0.00633408f
cc_302 N_MM7_g N_MS_1 0.00241719f
cc_303 N_MM7_g N_MS_11 0.00640431f
cc_304 N_MH_16 N_MS_18 0.00500454f
cc_305 N_MH_18 N_MS_14 0.00532125f
cc_306 N_MM7_g N_MM11_g 0.0293822f
x_PM_SDFHx1_ASAP7_75t_R%noxref_27 VSS N_noxref_27_1
+ PM_SDFHx1_ASAP7_75t_R%noxref_27
cc_307 N_noxref_27_1 N_MM22_g 0.00353394f
cc_308 N_noxref_27_1 N_CLKB_20 0.000167771f
cc_309 N_noxref_27_1 N_CLKB_7 0.000440498f
cc_310 N_noxref_27_1 N_CLKB_19 0.0269828f
cc_311 N_noxref_27_1 N_NET0120_8 0.000588553f
cc_312 N_noxref_27_1 N_noxref_26_1 0.00148613f
x_PM_SDFHx1_ASAP7_75t_R%noxref_29 VSS N_noxref_29_1
+ PM_SDFHx1_ASAP7_75t_R%noxref_29
cc_313 N_noxref_29_1 N_MM3_g 0.00150426f
cc_314 N_noxref_29_1 N_CLKB_7 0.000102268f
cc_315 N_noxref_29_1 N_CLKB_19 0.000579801f
cc_316 N_noxref_29_1 N_NET0120_8 0.0360113f
cc_317 N_noxref_29_1 N_noxref_26_1 0.000466399f
cc_318 N_noxref_29_1 N_noxref_27_1 0.00771781f
cc_319 N_noxref_29_1 N_noxref_28_1 0.00123926f
x_PM_SDFHx1_ASAP7_75t_R%noxref_30 VSS N_noxref_30_1
+ PM_SDFHx1_ASAP7_75t_R%noxref_30
cc_320 N_noxref_30_1 N_MM27_g 0.00149576f
cc_321 N_noxref_30_1 N_SI_1 0.00245483f
cc_322 N_noxref_30_1 N_CLKB_1 0.000184853f
cc_323 N_noxref_30_1 N_MM1_g 0.0107825f
cc_324 N_noxref_30_1 N_NET0120_2 0.0011575f
cc_325 N_noxref_30_1 N_NET0120_10 0.0161624f
cc_326 N_noxref_30_1 N_NET0120_9 0.0552254f
cc_327 N_noxref_30_1 N_NET0167_8 0.0371005f
x_PM_SDFHx1_ASAP7_75t_R%NET0118 VSS N_MM29_d N_MM5_d N_MM4_s N_NET0118_8
+ N_NET0118_9 N_NET0118_2 N_NET0118_7 N_NET0118_1 PM_SDFHx1_ASAP7_75t_R%NET0118
cc_328 N_NET0118_8 N_CLKN_2 0.000900373f
cc_329 N_NET0118_9 N_CLKN_25 0.000624583f
cc_330 N_NET0118_9 N_CLKN_20 0.000736306f
cc_331 N_NET0118_2 N_MM10_g 0.000868263f
cc_332 N_NET0118_8 N_MM10_g 0.0328318f
cc_333 N_NET0118_9 N_SE_13 0.00225598f
cc_334 N_NET0118_9 N_MM2_g 0.000313116f
cc_335 N_NET0118_9 N_SEN_14 0.000702422f
cc_336 N_NET0118_9 N_SEN_16 0.00364527f
cc_337 N_NET0118_9 N_D_4 0.000750205f
cc_338 N_NET0118_9 N_D_5 0.000763703f
cc_339 N_NET0118_7 N_D_1 0.000894976f
cc_340 N_NET0118_1 N_MM26_g 0.0011756f
cc_341 N_NET0118_7 N_MM26_g 0.0343743f
cc_342 N_NET0118_9 N_SI_4 0.000469266f
cc_343 N_NET0118_1 N_MM27_g 0.000780529f
cc_344 N_NET0118_7 N_SI_1 0.000842125f
cc_345 N_NET0118_9 N_SI_7 0.00284602f
cc_346 N_NET0118_7 N_MM27_g 0.0341056f
cc_347 N_NET0118_8 N_CLKB_21 0.000153102f
cc_348 N_NET0118_8 N_CLKB_1 0.0011175f
cc_349 N_NET0118_2 N_MM1_g 0.00116991f
cc_350 N_NET0118_9 N_CLKB_21 0.00228646f
cc_351 N_NET0118_8 N_MM1_g 0.0356602f
cc_352 N_NET0118_8 N_MH_10 0.0011512f
cc_353 N_NET0118_9 N_MH_15 0.000938035f
cc_354 N_NET0118_2 N_MH_4 0.00369322f
cc_355 N_NET0118_7 N_NET0167_8 0.000644414f
cc_356 N_NET0118_1 N_NET0167_10 0.000681134f
cc_357 N_NET0118_1 N_NET0167_2 0.00383264f
cc_358 N_NET0118_9 N_NET0167_10 0.00985153f
x_PM_SDFHx1_ASAP7_75t_R%SE VSS SE N_MM3_g N_MM30_g N_SE_11 N_SE_10 N_SE_7
+ N_SE_13 N_SE_8 N_SE_9 N_SE_12 N_SE_2 N_SE_1 PM_SDFHx1_ASAP7_75t_R%SE
cc_359 N_SE_11 N_CLKN_1 3.66328e-20
cc_360 N_SE_10 N_CLKN_22 4.43168e-20
cc_361 N_SE_11 N_CLKN_19 4.62706e-20
cc_362 N_SE_11 N_CLKN_18 5.29021e-20
cc_363 N_SE_7 N_CLKN_25 0.000377333f
cc_364 N_SE_11 N_CLKN_25 0.0003084f
cc_365 N_SE_13 N_CLKN_21 0.000482933f
cc_366 N_SE_13 N_CLKN_25 0.00183052f
cc_367 N_SE_8 N_CLKN_25 0.00288856f
x_PM_SDFHx1_ASAP7_75t_R%SH VSS N_MM14_g N_MM24_g N_MM13_s N_MM18_d N_MM12_s
+ N_MM17_d N_SH_6 N_SH_13 N_SH_14 N_SH_21 N_SH_15 N_SH_23 N_SH_17 N_SH_16
+ N_SH_5 N_SH_25 N_SH_20 N_SH_2 N_SH_22 N_SH_1 N_SH_18 N_SH_19 N_SH_24
+ PM_SDFHx1_ASAP7_75t_R%SH
cc_368 N_SH_6 N_MM17_g 0.000158318f
cc_369 N_SH_13 N_MM17_g 0.00676966f
cc_370 N_SH_14 N_MM17_g 0.00683991f
cc_371 N_SH_21 N_CLKN_21 0.000283052f
cc_372 N_SH_15 N_CLKN_21 0.000369575f
cc_373 N_SH_23 N_CLKN_21 0.000402567f
cc_374 N_SH_17 N_CLKN_21 0.000461538f
cc_375 N_SH_16 N_CLKN_3 0.000570191f
cc_376 N_SH_5 N_CLKN_3 0.000576027f
cc_377 N_SH_25 N_CLKN_25 0.000766503f
cc_378 N_SH_15 N_CLKN_25 0.00104611f
cc_379 N_SH_16 N_CLKN_21 0.00456887f
cc_380 N_SH_5 N_MM17_g 0.0183284f
cc_381 N_SH_20 N_SE_12 0.000222728f
cc_382 N_SH_16 N_SE_13 0.000315749f
cc_383 N_SH_2 N_SE_2 0.00163336f
cc_384 N_SH_15 N_SE_13 0.00103284f
cc_385 N_SH_25 N_SE_13 0.00207146f
cc_386 N_SH_22 N_SE_13 0.00268812f
cc_387 N_MM24_g N_MM30_g 0.00334156f
cc_388 N_SH_20 N_SE_9 0.0060972f
cc_389 N_SH_16 N_SEN_13 6.26363e-20
cc_390 N_MM24_g N_SEN_3 6.71442e-20
cc_391 N_SH_1 N_SEN_13 8.2894e-20
cc_392 N_SH_18 N_SEN_16 0.000109197f
cc_393 N_SH_25 N_SEN_15 0.000118258f
cc_394 N_SH_20 N_SEN_13 0.000157164f
cc_395 N_SH_25 N_SEN_13 0.00156706f
cc_396 N_SH_20 N_SEN_15 0.000255998f
cc_397 N_SH_19 N_SEN_16 0.000283404f
cc_398 N_SH_15 N_SEN_16 0.000374541f
cc_399 N_SH_25 N_SEN_16 0.00455622f
cc_400 N_SH_16 N_SEN_16 0.00610989f
cc_401 N_SH_14 N_CLKB_8 8.59205e-20
cc_402 N_SH_15 N_CLKB_26 8.92718e-20
cc_403 N_SH_21 N_CLKB_8 0.000196878f
cc_404 N_SH_23 N_CLKB_8 0.000203975f
cc_405 N_SH_13 N_MM12_g 0.00680288f
cc_406 N_SH_6 N_CLKB_8 0.000276286f
cc_407 N_SH_18 N_CLKB_8 0.000396208f
cc_408 N_SH_16 N_CLKB_8 0.000448364f
cc_409 N_SH_17 N_CLKB_8 0.00059347f
cc_410 N_SH_14 N_CLKB_4 0.000673075f
cc_411 N_SH_6 N_MM18_g 0.00100239f
cc_412 N_SH_5 N_CLKB_8 0.00282992f
cc_413 N_SH_5 N_MM12_g 0.00947788f
cc_414 N_SH_14 N_MM18_g 0.016093f
cc_415 N_SH_21 N_MS_3 0.00017983f
cc_416 N_SH_14 N_MS_3 0.000436412f
cc_417 N_SH_6 N_MS_3 0.000220843f
cc_418 N_SH_13 N_MS_3 0.000232021f
cc_419 N_SH_13 N_MS_11 0.000234021f
cc_420 N_SH_21 N_MS_4 0.000335704f
cc_421 N_SH_6 N_MS_4 0.000424812f
cc_422 N_SH_15 N_MS_16 0.000438227f
cc_423 N_SH_21 N_MS_17 0.00054066f
cc_424 N_SH_14 N_MS_4 0.000593146f
cc_425 N_SH_15 N_MS_19 0.00132359f
cc_426 N_SH_5 N_MS_3 0.00381434f
cc_427 N_SH_17 N_MM16_g 9.92271e-20
cc_428 N_SH_19 N_SS_13 0.000311072f
cc_429 N_MM14_g N_SS_3 0.000322929f
cc_430 N_MM14_g N_SS_4 0.00042065f
cc_431 N_SH_22 N_SS_15 0.000580125f
cc_432 N_SH_24 N_SS_16 0.000641453f
cc_433 N_SH_24 N_SS_14 0.00069774f
cc_434 N_SH_16 N_SS_1 0.000810777f
cc_435 N_SH_1 N_SS_14 0.000948913f
cc_436 N_MM14_g N_SS_1 0.00111318f
cc_437 N_SH_1 N_MM16_g 0.00135492f
cc_438 N_SH_18 N_SS_12 0.00154855f
cc_439 N_SH_25 N_SS_14 0.00175086f
cc_440 N_MM14_g N_SS_10 0.00649587f
cc_441 N_MM14_g N_SS_11 0.00660051f
cc_442 N_SH_16 N_SS_12 0.00462671f
cc_443 N_SH_19 N_SS_14 0.00483166f
cc_444 N_MM14_g N_MM16_g 0.0300176f
x_PM_SDFHx1_ASAP7_75t_R%CLKB VSS N_MM1_g N_MM9_g N_MM12_g N_MM18_g N_MM23_d
+ N_MM22_d N_CLKB_19 N_CLKB_20 N_CLKB_18 N_CLKB_26 N_CLKB_7 N_CLKB_6 N_CLKB_23
+ N_CLKB_24 N_CLKB_4 N_CLKB_22 N_CLKB_21 N_CLKB_8 N_CLKB_2 N_CLKB_1 N_CLKB_25
+ PM_SDFHx1_ASAP7_75t_R%CLKB
cc_445 N_CLKB_19 N_CLK_8 6.5469e-20
cc_446 N_CLKB_20 N_CLK_8 0.000230667f
cc_447 N_CLKB_18 N_CLK_8 8.77923e-20
cc_448 N_CLKB_26 N_CLK_8 0.000104577f
cc_449 N_CLKB_7 N_CLK_8 0.000350971f
cc_450 N_CLKB_6 N_CLK_8 0.000386451f
cc_451 N_CLKB_23 N_CLK_8 0.000352531f
cc_452 N_CLKB_20 N_CLK_6 0.000495512f
cc_453 N_CLKB_23 N_CLK_5 0.00140612f
cc_454 N_CLKB_24 N_CLK_8 0.00173679f
cc_455 N_CLKB_6 N_CLKN_25 5.40376e-20
cc_456 N_CLKB_7 N_MM22_g 0.000726602f
cc_457 N_CLKB_7 N_CLKN_18 8.53713e-20
cc_458 N_CLKB_4 N_MM17_g 0.000208159f
cc_459 N_CLKB_22 N_CLKN_25 0.000605602f
cc_460 N_CLKB_23 N_CLKN_19 0.000296518f
cc_461 N_CLKB_24 N_CLKN_19 0.000298484f
cc_462 N_CLKB_21 N_CLKN_25 0.000320154f
cc_463 N_CLKB_20 N_CLKN_19 0.0045855f
cc_464 N_CLKB_18 N_MM22_g 0.038648f
cc_465 N_CLKB_19 N_MM22_g 0.0111472f
cc_466 N_CLKB_26 N_CLKN_20 0.000466133f
cc_467 N_CLKB_8 N_CLKN_21 0.000531969f
cc_468 N_CLKB_20 N_CLKN_25 0.000540592f
cc_469 N_CLKB_2 N_MM10_g 0.000560135f
cc_470 N_CLKB_6 N_MM22_g 0.000598193f
cc_471 N_CLKB_20 N_CLKN_1 0.000615841f
cc_472 N_CLKB_8 N_CLKN_3 0.0027913f
cc_473 N_CLKB_19 N_CLKN_1 0.000777956f
cc_474 N_CLKB_1 N_CLKN_2 0.0022202f
cc_475 N_CLKB_25 N_CLKN_24 0.00165435f
cc_476 N_CLKB_21 N_CLKN_20 0.00255843f
cc_477 N_MM9_g N_MM10_g 0.00370396f
cc_478 N_CLKB_8 N_MM17_g 0.00493034f
cc_479 N_MM18_g N_MM17_g 0.00578926f
cc_480 N_MM1_g N_MM10_g 0.00704634f
cc_481 N_MM12_g N_MM17_g 0.0182757f
cc_482 N_CLKB_26 N_CLKN_25 0.0453372f
cc_483 N_CLKB_7 N_SE_11 5.05797e-20
cc_484 N_CLKB_6 N_SE_10 5.44239e-20
cc_485 N_MM18_g N_SE_13 0.000105906f
cc_486 N_CLKB_6 N_SE_7 0.000174715f
cc_487 N_CLKB_26 N_SE_13 0.000257394f
cc_488 N_CLKB_20 N_SE_7 0.0029933f
cc_489 N_CLKB_21 N_SE_13 0.000783418f
cc_490 N_CLKB_26 N_SE_8 0.00115164f
cc_491 N_CLKB_23 N_SE_10 0.00175627f
cc_492 N_CLKB_20 N_SE_11 0.00631258f
cc_493 N_MM1_g N_SI_5 7.69082e-20
cc_494 N_CLKB_1 N_SI_5 0.000397211f
cc_495 N_CLKB_26 N_SI_4 0.000310552f
cc_496 N_CLKB_26 N_SI_6 0.000321446f
cc_497 N_CLKB_21 N_SI_8 0.000647515f
cc_498 N_CLKB_21 N_SI_7 0.00068986f
cc_499 N_CLKB_25 N_SI_6 0.000925342f
cc_500 N_CLKB_26 N_SI_8 0.000957281f
cc_501 N_CLKB_21 N_SI_5 0.00302783f
*END of SDFHx1_ASAP7_75t_R.pxi
.ENDS
** Design:	SDFHx2_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "SDFHx2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "SDFHx2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_SDFHx2_ASAP7_75t_R%NET0167 VSS 2 3 1
c1 1 VSS 0.000995612f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3780 $Y2=0.0675
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%D VSS 4 3 1 5
c1 1 VSS 0.00721416f
c2 3 VSS 0.0461982f
c3 4 VSS 0.00468114f
c4 5 VSS 0.00360357f
r1 5 7 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.1080 $X2=0.4050 $Y2=0.1215
r2 4 7 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1215
r3 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r4 4 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%NET0166 VSS 14 27 7 9 1 11 12 10 8 2
c1 1 VSS 0.00638383f
c2 2 VSS 0.00557169f
c3 7 VSS 0.00466765f
c4 8 VSS 0.00320406f
c5 9 VSS 0.000876872f
c6 10 VSS 0.0175283f
c7 11 VSS 0.00129855f
c8 12 VSS 0.0020726f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0675 $X2=0.4840 $Y2=0.0675
r2 27 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4715 $Y2=0.0675
r3 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0675
+ $X2=0.4860 $Y2=0.0360
r4 23 24 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4475
+ $Y=0.0360 $X2=0.4860 $Y2=0.0360
r5 22 23 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4070
+ $Y=0.0360 $X2=0.4475 $Y2=0.0360
r6 21 22 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.3875
+ $Y=0.0360 $X2=0.4070 $Y2=0.0360
r7 20 21 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3605
+ $Y=0.0360 $X2=0.3875 $Y2=0.0360
r8 19 20 7.92845 $w=1.3e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3265
+ $Y=0.0360 $X2=0.3605 $Y2=0.0360
r9 10 12 1.03257 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3085 $Y=0.0360 $X2=0.2970 $Y2=0.0360
r10 10 19 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3085
+ $Y=0.0360 $X2=0.3265 $Y2=0.0360
r11 12 18 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.2970 $Y2=0.0540
r12 9 17 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0720 $X2=0.2970 $Y2=0.0900
r13 9 18 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0720 $X2=0.2970 $Y2=0.0540
r14 16 17 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2835 $Y=0.0900 $X2=0.2970 $Y2=0.0900
r15 11 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0900 $X2=0.2835 $Y2=0.0900
r16 11 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0900
+ $X2=0.2700 $Y2=0.0945
r17 1 15 23.8708 $w=2.02e-08 $l=4.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.2700 $Y=0.0540 $X2=0.2700 $Y2=0.0945
r18 14 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r19 7 13 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r20 1 7 1e-05
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%noxref_33 VSS 1
c1 1 VSS 0.00362774f
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%noxref_34 VSS 1
c1 1 VSS 0.00398969f
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.00420909f
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.00426895f
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%PD4 VSS 2 4 1
c1 1 VSS 0.00102981f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9890 $Y=0.2295 $X2=0.9765 $Y2=0.2295
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9550 $Y=0.2295 $X2=0.9595 $Y2=0.2295
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9595 $Y=0.2295 $X2=0.9765 $Y2=0.2295
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%PD3 VSS 2 4 1
c1 1 VSS 0.000910322f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.0405 $X2=0.7065 $Y2=0.0405
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.0405 $X2=0.6895 $Y2=0.0405
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6895 $Y=0.0405 $X2=0.7065 $Y2=0.0405
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%CLK VSS 13 3 4 6 1 5
c1 1 VSS 0.00302333f
c2 3 VSS 0.0599444f
c3 4 VSS 0.00256042f
c4 5 VSS 0.00482932f
c5 6 VSS 0.00193546f
r1 5 16 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0630 $X2=0.1080 $Y2=0.0900
r2 15 16 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.0900 $X2=0.1080 $Y2=0.0900
r3 6 9 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0900 $X2=0.0810 $Y2=0.1100
r4 6 15 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0900 $X2=0.0945 $Y2=0.0900
r5 13 12 2.73998 $w=1.3e-08 $l=1.18e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1900 $X2=0.0810 $Y2=0.1782
r6 11 12 3.20636 $w=1.3e-08 $l=1.37e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1645 $X2=0.0810 $Y2=0.1782
r7 10 11 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1530 $X2=0.0810 $Y2=0.1645
r8 8 10 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1530
r9 4 8 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1235 $X2=0.0810 $Y2=0.1350
r10 4 9 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1235 $X2=0.0810 $Y2=0.1100
r11 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r12 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%SI VSS 14 3 5 1 4 6 7
c1 1 VSS 0.00580989f
c2 3 VSS 0.00732761f
c3 4 VSS 0.00311399f
c4 5 VSS 0.00301514f
c5 6 VSS 0.00357509f
c6 7 VSS 0.00367721f
r1 6 19 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1980 $X2=0.5130 $Y2=0.1765
r2 5 7 3.2503 $w=1.53684e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1540 $X2=0.5130 $Y2=0.1350
r3 5 19 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1540 $X2=0.5130 $Y2=0.1765
r4 7 16 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1350 $X2=0.4945 $Y2=0.1350
r5 15 16 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4845
+ $Y=0.1350 $X2=0.4945 $Y2=0.1350
r6 14 15 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4750
+ $Y=0.1350 $X2=0.4845 $Y2=0.1350
r7 14 4 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4750
+ $Y=0.1350 $X2=0.4635 $Y2=0.1350
r8 14 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4750 $Y=0.1350
+ $X2=0.4790 $Y2=0.1350
r9 11 12 4.43042 $w=1.53e-08 $l=7.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.4715
+ $Y=0.1350 $X2=0.4790 $Y2=0.1350
r10 9 11 1.86855 $w=1.78125e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.4675 $Y=0.1350 $X2=0.4715 $Y2=0.1350
r11 1 9 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.4575
+ $Y=0.1350 $X2=0.4675 $Y2=0.1350
r12 3 1 2.53453 $w=1.32811e-07 $l=1.5e-09 $layer=LIG $thickness=5.23243e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4575 $Y2=0.1350
r13 3 11 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4715 $Y2=0.1350
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%noxref_26 VSS 1
c1 1 VSS 0.00433727f
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%noxref_28 VSS 1
c1 1 VSS 0.00582527f
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%noxref_29 VSS 1
c1 1 VSS 0.00587615f
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%noxref_30 VSS 1
c1 1 VSS 0.0126273f
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%PD2 VSS 7 12 4 5 1
c1 1 VSS 0.00742682f
c2 4 VSS 0.00184303f
c3 5 VSS 0.00234084f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7040 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r3 9 5 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.6765
+ $Y=0.2295 $X2=0.7020 $Y2=0.2295
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.6615
+ $Y=0.2295 $X2=0.6765 $Y2=0.2295
r5 1 8 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.6480
+ $Y=0.2295 $X2=0.6615 $Y2=0.2295
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.2295 $X2=0.6460 $Y2=0.2295
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.2295 $X2=0.6335 $Y2=0.2295
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%MH VSS 9 55 59 62 66 10 20 14 12 16 3 4 18 17 21
+ 1 19 15
c1 1 VSS 0.000217926f
c2 3 VSS 0.00474243f
c3 4 VSS 0.00496641f
c4 9 VSS 0.0361784f
c5 10 VSS 0.00228149f
c6 11 VSS 0.000103851f
c7 12 VSS 0.00212182f
c8 13 VSS 7.10038e-20
c9 14 VSS 0.00938877f
c10 15 VSS 0.00777006f
c11 16 VSS 0.00174916f
c12 17 VSS 0.000662745f
c13 18 VSS 0.000937044f
c14 19 VSS 0.00298925f
c15 20 VSS 5.96173e-20
c16 21 VSS 0.002694f
r1 66 65 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.2295 $X2=0.6085 $Y2=0.2295
r2 64 65 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6040 $Y=0.2295 $X2=0.6085 $Y2=0.2295
r3 3 64 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5920 $Y=0.2295 $X2=0.6040 $Y2=0.2295
r4 13 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2295 $X2=0.5920 $Y2=0.2295
r5 60 61 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.1890 $X2=0.5840 $Y2=0.1890
r6 62 60 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.1890 $X2=0.5795 $Y2=0.1890
r7 12 61 0.185185 $w=5.4e-08 $l=1e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.1890 $X2=0.5840 $Y2=0.1890
r8 12 3 0.518519 $w=3.9e-08 $l=4.05494e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.1890 $X2=0.5920 $Y2=0.2295
r9 59 58 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r10 57 58 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6580 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r11 4 57 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6460 $Y=0.0405 $X2=0.6580 $Y2=0.0405
r12 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0405 $X2=0.6460 $Y2=0.0405
r13 10 4 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0810 $X2=0.6460 $Y2=0.0810
r14 55 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.0810 $X2=0.6335 $Y2=0.0810
r15 3 47 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2295
+ $X2=0.5900 $Y2=0.2340
r16 4 41 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.0405
+ $X2=0.6440 $Y2=0.0360
r17 44 45 1.63233 $w=1.3e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.5990
+ $Y=0.2340 $X2=0.6060 $Y2=0.2340
r18 44 47 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5990
+ $Y=0.2340 $X2=0.5900 $Y2=0.2340
r19 43 45 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.6105
+ $Y=0.2340 $X2=0.6060 $Y2=0.2340
r20 42 43 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6305
+ $Y=0.2340 $X2=0.6105 $Y2=0.2340
r21 14 21 4.53042 $w=1.46981e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6665 $Y=0.2340 $X2=0.6930 $Y2=0.2340
r22 14 42 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.6665
+ $Y=0.2340 $X2=0.6305 $Y2=0.2340
r23 15 39 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.6530
+ $Y=0.0360 $X2=0.6705 $Y2=0.0360
r24 15 41 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6530
+ $Y=0.0360 $X2=0.6440 $Y2=0.0360
r25 21 38 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.2340 $X2=0.6930 $Y2=0.2160
r26 19 33 2.43171 $w=1.804e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6930 $Y=0.0360 $X2=0.6930 $Y2=0.0535
r27 19 39 3.59766 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.0360 $X2=0.6705 $Y2=0.0360
r28 37 38 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1980 $X2=0.6930 $Y2=0.2160
r29 36 37 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1800 $X2=0.6930 $Y2=0.1980
r30 35 36 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1680 $X2=0.6930 $Y2=0.1800
r31 34 35 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1590 $X2=0.6930 $Y2=0.1680
r32 17 20 2.43413 $w=1.59032e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6930 $Y=0.1465 $X2=0.6930 $Y2=0.1310
r33 17 34 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1465 $X2=0.6930 $Y2=0.1590
r34 32 33 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.0625 $X2=0.6930 $Y2=0.0535
r35 31 32 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.0720 $X2=0.6930 $Y2=0.0625
r36 30 31 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.0900 $X2=0.6930 $Y2=0.0720
r37 29 30 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1025 $X2=0.6930 $Y2=0.0900
r38 16 20 2.78392 $w=1.56471e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6930 $Y=0.1140 $X2=0.6930 $Y2=0.1310
r39 16 29 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1140 $X2=0.6930 $Y2=0.1025
r40 20 28 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1310 $X2=0.7110 $Y2=0.1310
r41 27 28 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1310 $X2=0.7110 $Y2=0.1310
r42 18 26 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.1310 $X2=0.7830 $Y2=0.1310
r43 18 27 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.1310 $X2=0.7290 $Y2=0.1310
r44 1 23 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.7830
+ $Y=0.1310 $X2=0.7830 $Y2=0.1310
r45 1 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7830 $Y=0.1310
+ $X2=0.7830 $Y2=0.1310
r46 9 23 0.314665 $w=2.27e-07 $l=4e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.7830 $Y=0.1350 $X2=0.7830 $Y2=0.1310
r47 3 12 1e-05
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%noxref_27 VSS 1
c1 1 VSS 0.00429947f
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%NET0141 VSS 12 13 27 28 7 9 1 2 8
c1 1 VSS 0.00532168f
c2 2 VSS 0.00532741f
c3 7 VSS 0.00334279f
c4 8 VSS 0.00336549f
c5 9 VSS 0.00269317f
r1 28 26 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r2 2 26 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r4 27 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r5 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4280 $Y2=0.1980
r6 21 22 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4185
+ $Y=0.1980 $X2=0.4280 $Y2=0.1980
r7 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1980 $X2=0.4185 $Y2=0.1980
r8 19 20 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.3875
+ $Y=0.1980 $X2=0.4050 $Y2=0.1980
r9 18 19 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3695
+ $Y=0.1980 $X2=0.3875 $Y2=0.1980
r10 17 18 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1980 $X2=0.3695 $Y2=0.1980
r11 16 17 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.1980 $X2=0.3510 $Y2=0.1980
r12 15 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1980 $X2=0.3375 $Y2=0.1980
r13 14 15 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3130
+ $Y=0.1980 $X2=0.3240 $Y2=0.1980
r14 9 14 0.699569 $w=1.3e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.3100
+ $Y=0.1980 $X2=0.3130 $Y2=0.1980
r15 1 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.1980
r16 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r17 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r18 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r19 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%MS VSS 10 43 46 50 52 13 17 19 18 3 15 12 1 11 4
+ 14 16
c1 1 VSS 0.00317511f
c2 3 VSS 0.00574969f
c3 4 VSS 0.00955833f
c4 10 VSS 0.0376963f
c5 11 VSS 0.00328742f
c6 12 VSS 0.00311932f
c7 13 VSS 0.00262986f
c8 14 VSS 0.000855738f
c9 15 VSS 0.00355241f
c10 16 VSS 0.00188609f
c11 17 VSS 0.00112546f
c12 18 VSS 0.00137227f
c13 19 VSS 0.00118266f
c14 20 VSS 0.00294898f
r1 52 51 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8810 $Y=0.2295 $X2=0.8785 $Y2=0.2295
r2 13 51 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8660 $Y=0.2295 $X2=0.8785 $Y2=0.2295
r3 12 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.2295 $X2=0.8080 $Y2=0.2295
r4 50 12 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.2295 $X2=0.7955 $Y2=0.2295
r5 47 13 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8370 $Y=0.2295 $X2=0.8640 $Y2=0.2295
r6 4 47 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08 $X=0.8100
+ $Y=0.2295 $X2=0.8370 $Y2=0.2295
r7 4 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8100 $Y=0.2295
+ $X2=0.8100 $Y2=0.2340
r8 15 20 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.2340 $X2=0.8370 $Y2=0.2340
r9 46 45 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8270 $Y=0.0405 $X2=0.8245 $Y2=0.0405
r10 44 45 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8200 $Y=0.0405 $X2=0.8245 $Y2=0.0405
r11 3 44 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8080 $Y=0.0405 $X2=0.8200 $Y2=0.0405
r12 11 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.0405 $X2=0.8080 $Y2=0.0405
r13 43 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.0405 $X2=0.7955 $Y2=0.0405
r14 20 39 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.2340 $X2=0.8370 $Y2=0.2160
r15 3 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8100 $Y=0.0405
+ $X2=0.8100 $Y2=0.0535
r16 38 39 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1870 $X2=0.8370 $Y2=0.2160
r17 37 38 4.89699 $w=1.3e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1660 $X2=0.8370 $Y2=0.1870
r18 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1525 $X2=0.8370 $Y2=0.1660
r19 35 36 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1310 $X2=0.8370 $Y2=0.1525
r20 34 35 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1115 $X2=0.8370 $Y2=0.1310
r21 17 31 1.15159 $w=1.75e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1000 $X2=0.8370 $Y2=0.0900
r22 17 34 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1000 $X2=0.8370 $Y2=0.1115
r23 16 32 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0625 $X2=0.8100 $Y2=0.0720
r24 16 33 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0625 $X2=0.8100 $Y2=0.0535
r25 30 31 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8235 $Y=0.0900 $X2=0.8370 $Y2=0.0900
r26 19 28 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.0900 $X2=0.7965 $Y2=0.0900
r27 19 30 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.0900 $X2=0.8235 $Y2=0.0900
r28 19 32 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0900 $X2=0.8100 $Y2=0.0720
r29 27 28 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.7740
+ $Y=0.0900 $X2=0.7965 $Y2=0.0900
r30 14 27 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7470
+ $Y=0.0900 $X2=0.7740 $Y2=0.0900
r31 14 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7470 $Y=0.0900
+ $X2=0.7500 $Y2=0.0900
r32 14 18 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7470
+ $Y=0.0900 $X2=0.7290 $Y2=0.0900
r33 25 26 5.02115 $w=1.53e-08 $l=8.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.7415 $Y=0.0900 $X2=0.7500 $Y2=0.0900
r34 23 25 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.7385 $Y=0.0900 $X2=0.7415 $Y2=0.0900
r35 1 23 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.7285
+ $Y=0.0900 $X2=0.7385 $Y2=0.0900
r36 1 22 2.48102 $w=2.2e-08 $l=5e-10 $layer=LIG $thickness=4.8e-08 $X=0.7285
+ $Y=0.0900 $X2=0.7290 $Y2=0.0900
r37 22 25 1.47681 $w=1.53e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7290 $Y=0.0900 $X2=0.7415 $Y2=0.0900
r38 10 22 0.314665 $w=2.27e-07 $l=4.5e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.7290 $Y=0.1350 $X2=0.7290 $Y2=0.0900
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%NET0120 VSS 13 24 26 8 1 2 9 11 10
c1 1 VSS 0.00560869f
c2 2 VSS 0.0086144f
c3 8 VSS 0.00327637f
c4 9 VSS 0.00234801f
c5 10 VSS 0.0021375f
c6 11 VSS 0.0229327f
r1 26 25 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r2 10 25 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5420 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r3 9 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4840 $Y2=0.2025
r4 24 9 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r5 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5130 $Y=0.2025
+ $X2=0.4900 $Y2=0.2340
r6 20 21 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4810
+ $Y=0.2340 $X2=0.4900 $Y2=0.2340
r7 19 20 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4690
+ $Y=0.2340 $X2=0.4810 $Y2=0.2340
r8 18 19 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4540
+ $Y=0.2340 $X2=0.4690 $Y2=0.2340
r9 17 18 17.7224 $w=1.3e-08 $l=7.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.4540 $Y2=0.2340
r10 16 17 19.5879 $w=1.3e-08 $l=8.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2940
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r11 15 16 5.59655 $w=1.3e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.2940 $Y2=0.2340
r12 11 15 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2580
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r13 8 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2160
+ $X2=0.2700 $Y2=0.2340
r14 1 8 23.8708 $w=2.02e-08 $l=4.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.2700 $Y=0.1755 $X2=0.2700 $Y2=0.2160
r15 13 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r16 8 12 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r17 2 10 1e-05
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%NET0118 VSS 12 13 29 8 9 2 7 1
c1 1 VSS 0.00351716f
c2 2 VSS 0.00380905f
c3 7 VSS 0.0029416f
c4 8 VSS 0.00227395f
c5 9 VSS 0.0024397f
r1 29 28 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.0675 $X2=0.6085 $Y2=0.0675
r2 27 28 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6040 $Y=0.0675 $X2=0.6085 $Y2=0.0675
r3 8 27 0.123457 $w=8.1e-08 $l=1e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.0675 $X2=0.6040 $Y2=0.0675
r4 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0675
+ $X2=0.5900 $Y2=0.0720
r5 23 24 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.5805
+ $Y=0.0720 $X2=0.5900 $Y2=0.0720
r6 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0720 $X2=0.5805 $Y2=0.0720
r7 21 22 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.0720 $X2=0.5670 $Y2=0.0720
r8 20 21 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0720 $X2=0.5400 $Y2=0.0720
r9 19 20 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5020
+ $Y=0.0720 $X2=0.5130 $Y2=0.0720
r10 18 19 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4805
+ $Y=0.0720 $X2=0.5020 $Y2=0.0720
r11 17 18 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.4540
+ $Y=0.0720 $X2=0.4805 $Y2=0.0720
r12 16 17 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4440
+ $Y=0.0720 $X2=0.4540 $Y2=0.0720
r13 15 16 1.63233 $w=1.3e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.4370
+ $Y=0.0720 $X2=0.4440 $Y2=0.0720
r14 14 15 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4280
+ $Y=0.0720 $X2=0.4370 $Y2=0.0720
r15 9 14 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4205
+ $Y=0.0720 $X2=0.4280 $Y2=0.0720
r16 1 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4280 $Y2=0.0720
r17 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r18 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r19 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0675 $X2=0.4320 $Y2=0.0675
r20 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4175 $Y2=0.0675
r21 2 8 1e-05
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%noxref_31 VSS 1
c1 1 VSS 0.0035965f
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%SEN VSS 9 45 47 16 12 13 4 10 11 14 3 1 15
c1 1 VSS 0.00392947f
c2 3 VSS 0.00880265f
c3 4 VSS 0.00686648f
c4 9 VSS 0.0815982f
c5 10 VSS 0.00434231f
c6 11 VSS 0.004695f
c7 12 VSS 0.00182409f
c8 13 VSS 0.00383941f
c9 14 VSS 0.00083748f
c10 15 VSS 0.00591828f
c11 16 VSS 0.0164786f
r1 47 46 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.2050 $Y=0.2295 $X2=1.2025 $Y2=0.2295
r2 11 46 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.1900 $Y=0.2295 $X2=1.2025 $Y2=0.2295
r3 4 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.1880 $Y=0.2295
+ $X2=1.1880 $Y2=0.2340
r4 45 44 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.2050 $Y=0.0405 $X2=1.2025 $Y2=0.0405
r5 10 44 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.1900 $Y=0.0405 $X2=1.2025 $Y2=0.0405
r6 41 42 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.1745
+ $Y=0.2340 $X2=1.1880 $Y2=0.2340
r7 15 37 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1610 $Y=0.2340 $X2=1.1610 $Y2=0.2125
r8 15 41 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1610 $Y=0.2340 $X2=1.1745 $Y2=0.2340
r9 39 10 3.98201 $w=3.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.1730 $Y=0.0455 $X2=1.1880 $Y2=0.0455
r10 38 39 3.18561 $w=3.32e-08 $l=1.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.1610 $Y=0.0455 $X2=1.1730 $Y2=0.0455
r11 3 38 3.31834 $w=3.32e-08 $l=1.25e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.1485 $Y=0.0455 $X2=1.1610 $Y2=0.0455
r12 36 37 15.7403 $w=1.3e-08 $l=6.75e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.1450 $X2=1.1610 $Y2=0.2125
r13 35 36 14.9241 $w=1.3e-08 $l=6.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0810 $X2=1.1610 $Y2=0.1450
r14 34 35 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0650 $X2=1.1610 $Y2=0.0810
r15 33 34 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0515 $X2=1.1610 $Y2=0.0650
r16 33 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.1610 $Y=0.0515
+ $X2=1.1610 $Y2=0.0455
r17 32 33 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0425 $X2=1.1610 $Y2=0.0515
r18 13 32 1.28254 $w=1.3e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0370 $X2=1.1610 $Y2=0.0425
r19 30 35 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=1.1610 $Y=0.0810
+ $X2=1.1610 $Y2=0.0810
r20 29 30 27.2832 $w=1.3e-08 $l=1.17e-07 $layer=M2 $thickness=3.6e-08 $X=1.0440
+ $Y=0.0810 $X2=1.1610 $Y2=0.0810
r21 28 29 29.3819 $w=1.3e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.9180
+ $Y=0.0810 $X2=1.0440 $Y2=0.0810
r22 27 28 67.1587 $w=1.3e-08 $l=2.88e-07 $layer=M2 $thickness=3.6e-08 $X=0.6300
+ $Y=0.0810 $X2=0.9180 $Y2=0.0810
r23 26 27 65.0599 $w=1.3e-08 $l=2.79e-07 $layer=M2 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0810 $X2=0.6300 $Y2=0.0810
r24 16 26 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.3395
+ $Y=0.0810 $X2=0.3510 $Y2=0.0810
r25 14 22 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.0720 $X2=0.3510 $Y2=0.0855
r26 14 26 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.3510 $Y=0.0720 $X2=0.3510
+ $Y2=0.0810
r27 22 23 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0855 $X2=0.3510 $Y2=0.0945
r28 22 26 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.3510 $Y=0.0855 $X2=0.3510
+ $Y2=0.0810
r29 21 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1080 $X2=0.3510 $Y2=0.0945
r30 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1215 $X2=0.3510 $Y2=0.1080
r31 12 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1215
r32 9 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r33 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
r34 4 11 1e-05
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%noxref_35 VSS 1
c1 1 VSS 0.0423882f
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%QN VSS 22 16 17 28 29 9 7 8 10 11 1 2
c1 1 VSS 0.0102161f
c2 2 VSS 0.0103336f
c3 7 VSS 0.00453286f
c4 8 VSS 0.00449267f
c5 9 VSS 0.00924125f
c6 10 VSS 0.00919134f
c7 11 VSS 0.00730058f
c8 12 VSS 0.00338762f
c9 13 VSS 0.00335107f
r1 29 27 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.3130 $Y=0.2025 $X2=1.3105 $Y2=0.2025
r2 2 27 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.2960 $Y=0.2025 $X2=1.3105 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.2815 $Y=0.2025 $X2=1.2960 $Y2=0.2025
r4 28 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.2790 $Y=0.2025 $X2=1.2815 $Y2=0.2025
r5 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.2960 $Y=0.2025
+ $X2=1.2960 $Y2=0.2340
r6 24 25 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=1.2960
+ $Y=0.2340 $X2=1.3365 $Y2=0.2340
r7 10 24 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.2845
+ $Y=0.2340 $X2=1.2960 $Y2=0.2340
r8 13 23 0.624487 $w=2.20462e-08 $l=9.8e-09 $layer=M1 $thickness=3.6e-08
+ $X=1.3770 $Y=0.2340 $X2=1.3770 $Y2=0.2242
r9 13 25 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3770 $Y=0.2340 $X2=1.3365 $Y2=0.2340
r10 22 23 0.291487 $w=1.3e-08 $l=1.2e-09 $layer=M1 $thickness=3.6e-08 $X=1.3770
+ $Y=0.2230 $X2=1.3770 $Y2=0.2242
r11 22 21 2.73998 $w=1.3e-08 $l=1.18e-08 $layer=M1 $thickness=3.6e-08 $X=1.3770
+ $Y=0.2230 $X2=1.3770 $Y2=0.2112
r12 20 21 15.4488 $w=1.3e-08 $l=6.62e-08 $layer=M1 $thickness=3.6e-08 $X=1.3770
+ $Y=0.1450 $X2=1.3770 $Y2=0.2112
r13 11 12 5.69636 $w=1.58e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3770 $Y=0.0675 $X2=1.3770 $Y2=0.0360
r14 11 20 18.0722 $w=1.3e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=1.3770
+ $Y=0.0675 $X2=1.3770 $Y2=0.1450
r15 12 19 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3770 $Y=0.0360 $X2=1.3365 $Y2=0.0360
r16 18 19 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=1.2960
+ $Y=0.0360 $X2=1.3365 $Y2=0.0360
r17 9 18 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.2845
+ $Y=0.0360 $X2=1.2960 $Y2=0.0360
r18 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.2960 $Y=0.0675
+ $X2=1.2960 $Y2=0.0360
r19 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.3130 $Y=0.0675 $X2=1.3105 $Y2=0.0675
r20 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.2960 $Y=0.0675 $X2=1.3105 $Y2=0.0675
r21 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.2815 $Y=0.0675 $X2=1.2960 $Y2=0.0675
r22 16 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.2790 $Y=0.0675 $X2=1.2815 $Y2=0.0675
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%noxref_36 VSS 1
c1 1 VSS 0.0423658f
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%PD5 VSS 7 12 4 1 5
c1 1 VSS 0.00742971f
c2 4 VSS 0.00187924f
c3 5 VSS 0.00237018f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9890 $Y=0.0405 $X2=0.9865 $Y2=0.0405
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9740 $Y=0.0405 $X2=0.9865 $Y2=0.0405
r3 9 5 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.9585
+ $Y=0.0405 $X2=0.9720 $Y2=0.0405
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.9435
+ $Y=0.0405 $X2=0.9585 $Y2=0.0405
r5 1 8 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.9180
+ $Y=0.0405 $X2=0.9435 $Y2=0.0405
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9035 $Y=0.0405 $X2=0.9160 $Y2=0.0405
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9010 $Y=0.0405 $X2=0.9035 $Y2=0.0405
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%noxref_32 VSS 1
c1 1 VSS 0.00379324f
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%CLKB VSS 14 15 16 17 85 87 26 19 7 18 24 6 20 23
+ 4 22 21 8 2 1 25
c1 1 VSS 0.000281941f
c2 2 VSS 6.4568e-20
c3 3 VSS 1e-36
c4 4 VSS 0.000306315f
c5 6 VSS 0.00736731f
c6 7 VSS 0.0074559f
c7 8 VSS 0.00383894f
c8 14 VSS 0.00583847f
c9 15 VSS 0.00508968f
c10 16 VSS 0.0043852f
c11 17 VSS 0.00520976f
c12 18 VSS 0.00760048f
c13 19 VSS 0.00754538f
c14 20 VSS 0.00332891f
c15 21 VSS 0.00180989f
c16 22 VSS 0.00141674f
c17 23 VSS 0.00609749f
c18 24 VSS 0.00603675f
c19 25 VSS 0.000615203f
c20 26 VSS 0.0234915f
r1 19 7 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1600 $Y2=0.2160
r2 87 19 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r3 18 6 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1600 $Y2=0.0540
r4 85 18 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r5 7 80 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r6 6 77 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r7 1 72 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1355
+ $X2=0.5670 $Y2=0.1350
r8 14 1 3.19489 $w=1.24e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1355
r9 80 81 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r10 24 68 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.1890 $Y2=0.2160
r11 24 81 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2340 $X2=0.1755 $Y2=0.2340
r12 77 78 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r13 23 64 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1890 $Y2=0.0630
r14 23 78 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1755 $Y2=0.0360
r15 25 69 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.1980 $X2=0.5670 $Y2=0.1845
r16 25 54 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.5670 $Y=0.1980 $X2=0.5670
+ $Y2=0.1890
r17 72 73 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1485
r18 70 73 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1620 $X2=0.5670 $Y2=0.1485
r19 21 69 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1755 $X2=0.5670 $Y2=0.1845
r20 21 70 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1755 $X2=0.5670 $Y2=0.1620
r21 67 68 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2035 $X2=0.1890 $Y2=0.2160
r22 66 67 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1990 $X2=0.1890 $Y2=0.2035
r23 65 66 1.28254 $w=1.3e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1935 $X2=0.1890 $Y2=0.1990
r24 63 64 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0900 $X2=0.1890 $Y2=0.0630
r25 62 63 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1100 $X2=0.1890 $Y2=0.0900
r26 61 62 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1325 $X2=0.1890 $Y2=0.1100
r27 60 61 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1540 $X2=0.1890 $Y2=0.1325
r28 59 60 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1655 $X2=0.1890 $Y2=0.1540
r29 58 65 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1845 $X2=0.1890 $Y2=0.1935
r30 20 58 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1735 $X2=0.1890 $Y2=0.1845
r31 20 59 1.86552 $w=1.3e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1735 $X2=0.1890 $Y2=0.1655
r32 55 56 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.6480
+ $Y=0.1890 $X2=0.7290 $Y2=0.1890
r33 54 55 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1890 $X2=0.6480 $Y2=0.1890
r34 54 69 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.5670 $Y=0.1890 $X2=0.5670
+ $Y2=0.1845
r35 53 54 44.0729 $w=1.3e-08 $l=1.89e-07 $layer=M2 $thickness=3.6e-08 $X=0.3780
+ $Y=0.1890 $X2=0.5670 $Y2=0.1890
r36 52 53 44.0729 $w=1.3e-08 $l=1.89e-07 $layer=M2 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1890 $X2=0.3780 $Y2=0.1890
r37 52 58 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1890 $Y=0.1890
+ $X2=0.1890 $Y2=0.1845
r38 26 52 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.1775
+ $Y=0.1890 $X2=0.1890 $Y2=0.1890
r39 4 49 2.78395 $w=2.4e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.9450
+ $Y=0.1780 $X2=0.9450 $Y2=0.1780
r40 17 4 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.9450 $Y=0.1350 $X2=0.9450 $Y2=0.1780
r41 2 42 2.78395 $w=2.4e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.6750
+ $Y=0.1780 $X2=0.6750 $Y2=0.1780
r42 15 2 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.6750 $Y=0.1350 $X2=0.6750 $Y2=0.1780
r43 50 56 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.7290 $Y=0.1845
+ $X2=0.7290 $Y2=0.1890
r44 22 50 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1680 $X2=0.7290 $Y2=0.1845
r45 48 49 6.83711 $w=2.22e-08 $l=1.5e-09 $layer=LISD $thickness=2.7e-08
+ $X=0.9435 $Y=0.1780 $X2=0.9450 $Y2=0.1780
r46 47 48 12.9145 $w=2.22e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9180 $Y=0.1780 $X2=0.9435 $Y2=0.1780
r47 46 47 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9045 $Y=0.1780 $X2=0.9180 $Y2=0.1780
r48 45 46 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8910 $Y=0.1780 $X2=0.9045 $Y2=0.1780
r49 44 45 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8775 $Y=0.1780 $X2=0.8910 $Y2=0.1780
r50 43 44 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8640 $Y=0.1780 $X2=0.8775 $Y2=0.1780
r51 41 42 12.9145 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6885 $Y=0.1780 $X2=0.6750 $Y2=0.1780
r52 40 41 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7155 $Y=0.1780 $X2=0.6885 $Y2=0.1780
r53 38 39 6.07743 $w=2.22e-08 $l=1.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7290 $Y=0.1780 $X2=0.7410 $Y2=0.1780
r54 38 50 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7290 $Y=0.1780
+ $X2=0.7290 $Y2=0.1845
r55 37 38 5.31775 $w=2.22e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7185 $Y=0.1780 $X2=0.7290 $Y2=0.1780
r56 37 40 1.51936 $w=2.22e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.7185
+ $Y=0.1780 $X2=0.7155 $Y2=0.1780
r57 36 39 4.55807 $w=2.22e-08 $l=9e-09 $layer=LISD $thickness=2.7e-08 $X=0.7500
+ $Y=0.1780 $X2=0.7410 $Y2=0.1780
r58 35 36 6.07743 $w=2.22e-08 $l=1.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7620 $Y=0.1780 $X2=0.7500 $Y2=0.1780
r59 34 35 4.05162 $w=2.22e-08 $l=8e-09 $layer=LISD $thickness=2.7e-08 $X=0.7700
+ $Y=0.1780 $X2=0.7620 $Y2=0.1780
r60 33 34 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7835 $Y=0.1780 $X2=0.7700 $Y2=0.1780
r61 32 33 6.58388 $w=2.22e-08 $l=1.3e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7965 $Y=0.1780 $X2=0.7835 $Y2=0.1780
r62 31 32 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8100 $Y=0.1780 $X2=0.7965 $Y2=0.1780
r63 8 31 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8370 $Y=0.1780 $X2=0.8100 $Y2=0.1780
r64 8 43 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8370 $Y=0.1780 $X2=0.8640 $Y2=0.1780
r65 3 30 2.78395 $w=2.4e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.8370
+ $Y=0.1780 $X2=0.8370 $Y2=0.1780
r66 3 8 10.3807 $w=2.30357e-08 $l=0 $layer=LISD $thickness=3.675e-08 $X=0.8370
+ $Y=0.1780 $X2=0.8370 $Y2=0.1780
r67 16 30 0.314665 $w=2.27e-07 $l=4.3e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.8370 $Y=0.1350 $X2=0.8370 $Y2=0.1780
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%SS VSS 9 34 39 14 13 12 17 16 3 4 15 1 10 11
c1 1 VSS 0.00111191f
c2 3 VSS 0.00569209f
c3 4 VSS 0.00656443f
c4 9 VSS 0.0384075f
c5 10 VSS 0.00327151f
c6 11 VSS 0.00332018f
c7 12 VSS 0.000996925f
c8 13 VSS 0.00845958f
c9 14 VSS 0.00183764f
c10 15 VSS 0.00251762f
c11 16 VSS 0.00670785f
c12 17 VSS 0.0023053f
r1 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0655 $Y=0.2295 $X2=1.0780 $Y2=0.2295
r2 39 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0630 $Y=0.2295 $X2=1.0655 $Y2=0.2295
r3 4 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0800 $Y=0.2295
+ $X2=1.0800 $Y2=0.2340
r4 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.0800
+ $Y=0.2340 $X2=1.0935 $Y2=0.2340
r5 16 32 7.21452 $w=1.425e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.2340 $X2=1.1070 $Y2=0.1980
r6 16 37 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1070 $Y=0.2340 $X2=1.0935 $Y2=0.2340
r7 10 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.0655 $Y=0.0405 $X2=1.0780 $Y2=0.0405
r8 34 10 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.0630 $Y=0.0405 $X2=1.0655 $Y2=0.0405
r9 31 32 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.1440 $X2=1.1070 $Y2=0.1980
r10 14 30 8.95608 $w=1.36627e-08 $l=4.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1070 $Y=0.0810 $X2=1.1070 $Y2=0.0395
r11 14 31 14.691 $w=1.3e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.0810 $X2=1.1070 $Y2=0.1440
r12 3 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0800 $Y=0.0405
+ $X2=1.0800 $Y2=0.0360
r13 17 29 1.40651 $w=1.51875e-08 $l=1.45774e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1070 $Y=0.0305 $X2=1.0935 $Y2=0.0360
r14 17 30 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.0305 $X2=1.1070 $Y2=0.0395
r15 28 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.0800
+ $Y=0.0360 $X2=1.0935 $Y2=0.0360
r16 27 28 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.0685
+ $Y=0.0360 $X2=1.0800 $Y2=0.0360
r17 26 27 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.0640
+ $Y=0.0360 $X2=1.0685 $Y2=0.0360
r18 25 26 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.0360 $X2=1.0640 $Y2=0.0360
r19 13 15 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0260 $Y=0.0360 $X2=0.9990 $Y2=0.0360
r20 13 25 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.0360 $X2=1.0530 $Y2=0.0360
r21 12 22 8.04505 $w=1.3e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.9990
+ $Y=0.0705 $X2=0.9990 $Y2=0.1050
r22 12 15 6.39593 $w=1.55565e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9990 $Y=0.0705 $X2=0.9990 $Y2=0.0360
r23 1 19 2.36633 $w=2.3e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.9990
+ $Y=0.1055 $X2=0.9990 $Y2=0.1055
r24 1 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.9990 $Y=0.1055
+ $X2=0.9990 $Y2=0.1050
r25 9 19 0.314665 $w=2.27e-07 $l=2.95e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.9990 $Y=0.1350 $X2=0.9990 $Y2=0.1055
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%SH VSS 11 12 13 76 79 81 84 6 14 15 22 16 24 18
+ 17 5 26 21 2 23 1 19 20 25
c1 1 VSS 0.000689258f
c2 2 VSS 0.0076319f
c3 5 VSS 0.00498967f
c4 6 VSS 0.00514577f
c5 11 VSS 0.0378177f
c6 12 VSS 0.0803989f
c7 13 VSS 0.0809766f
c8 14 VSS 0.00503391f
c9 15 VSS 0.0052013f
c10 16 VSS 0.00800642f
c11 17 VSS 0.000583398f
c12 18 VSS 0.00157536f
c13 19 VSS 0.00122249f
c14 20 VSS 0.000193154f
c15 21 VSS 0.00461722f
c16 22 VSS 0.00671959f
c17 23 VSS 0.0022087f
c18 24 VSS 0.000162363f
c19 25 VSS 0.000441033f
c20 26 VSS 0.0154624f
r1 84 83 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8810 $Y=0.0405 $X2=0.8785 $Y2=0.0405
r2 5 83 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8660 $Y=0.0405 $X2=0.8785 $Y2=0.0405
r3 80 5 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8540 $Y=0.0405 $X2=0.8660 $Y2=0.0405
r4 14 80 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.0405 $X2=0.8540 $Y2=0.0405
r5 81 14 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.0405 $X2=0.8495 $Y2=0.0405
r6 79 78 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9350 $Y=0.2295 $X2=0.9325 $Y2=0.2295
r7 77 78 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9280 $Y=0.2295 $X2=0.9325 $Y2=0.2295
r8 6 77 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9160 $Y=0.2295 $X2=0.9280 $Y2=0.2295
r9 15 6 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9035 $Y=0.2295 $X2=0.9160 $Y2=0.2295
r10 76 15 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9010 $Y=0.2295 $X2=0.9035 $Y2=0.2295
r11 13 68 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=1.3230
+ $Y=0.1350 $X2=1.3230 $Y2=0.1360
r12 12 60 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=1.2690 $Y=0.1350 $X2=1.2690 $Y2=0.1360
r13 5 58 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.0405
+ $X2=0.8640 $Y2=0.0360
r14 6 53 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.9180 $Y=0.2295
+ $X2=0.9180 $Y2=0.2340
r15 66 68 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.3105 $Y=0.1360 $X2=1.3230 $Y2=0.1360
r16 65 66 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.2960 $Y=0.1360 $X2=1.3105 $Y2=0.1360
r17 63 65 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.2815 $Y=0.1360 $X2=1.2960 $Y2=0.1360
r18 61 63 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=1.2785 $Y=0.1360 $X2=1.2815 $Y2=0.1360
r19 60 61 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=1.2690
+ $Y=0.1360 $X2=1.2785 $Y2=0.1360
r20 2 60 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=1.2595
+ $Y=0.1360 $X2=1.2690 $Y2=0.1360
r21 58 59 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.0360 $X2=0.8775 $Y2=0.0360
r22 56 59 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.0360 $X2=0.8775 $Y2=0.0360
r23 55 56 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.9020
+ $Y=0.0360 $X2=0.8910 $Y2=0.0360
r24 16 23 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.9200
+ $Y=0.0360 $X2=0.9450 $Y2=0.0360
r25 16 55 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.9200
+ $Y=0.0360 $X2=0.9020 $Y2=0.0360
r26 53 54 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.2340 $X2=0.9315 $Y2=0.2340
r27 22 54 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.2340 $X2=0.9315 $Y2=0.2340
r28 50 60 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.2690 $Y=0.1445
+ $X2=1.2690 $Y2=0.1360
r29 21 50 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.2690
+ $Y=0.1085 $X2=1.2690 $Y2=0.1445
r30 23 44 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.0360 $X2=0.9450 $Y2=0.0630
r31 18 39 6.50021 $w=1.33448e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.1980 $X2=0.9450 $Y2=0.1690
r32 18 22 7.21452 $w=1.425e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.1980 $X2=0.9450 $Y2=0.2340
r33 48 50 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=1.2690 $Y=0.1530
+ $X2=1.2690 $Y2=0.1445
r34 47 48 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=1.2445
+ $Y=0.1530 $X2=1.2690 $Y2=0.1530
r35 46 47 9.91056 $w=1.3e-08 $l=4.25e-08 $layer=M2 $thickness=3.6e-08 $X=1.2020
+ $Y=0.1530 $X2=1.2445 $Y2=0.1530
r36 45 46 32.0636 $w=1.3e-08 $l=1.375e-07 $layer=M2 $thickness=3.6e-08
+ $X=1.0645 $Y=0.1530 $X2=1.2020 $Y2=0.1530
r37 26 45 27.8662 $w=1.3e-08 $l=1.195e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.9450 $Y=0.1530 $X2=1.0645 $Y2=0.1530
r38 26 40 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.9450 $Y=0.1530 $X2=0.9450
+ $Y2=0.1485
r39 43 44 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.0900 $X2=0.9450 $Y2=0.0630
r40 42 43 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1000 $X2=0.9450 $Y2=0.0900
r41 41 42 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1100 $X2=0.9450 $Y2=0.1000
r42 17 40 3.96423 $w=1.3e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1315 $X2=0.9450 $Y2=0.1485
r43 17 41 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1315 $X2=0.9450 $Y2=0.1100
r44 38 39 0.4592 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1645 $X2=0.9450 $Y2=0.1690
r45 24 38 0.714311 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1575 $X2=0.9450 $Y2=0.1645
r46 24 40 1.50855 $w=1.55e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1575 $X2=0.9450 $Y2=0.1485
r47 24 26 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.9450 $Y=0.1575 $X2=0.9450
+ $Y2=0.1530
r48 37 39 4.4015 $w=1.35e-08 $l=2.78927e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9720 $Y=0.1620 $X2=0.9450 $Y2=0.1690
r49 36 37 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9990
+ $Y=0.1620 $X2=0.9720 $Y2=0.1620
r50 19 25 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0260 $Y=0.1620 $X2=1.0530 $Y2=0.1620
r51 19 36 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.1620 $X2=0.9990 $Y2=0.1620
r52 25 34 0.915974 $w=2.10182e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0530 $Y=0.1620 $X2=1.0530 $Y2=0.1510
r53 33 34 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1400 $X2=1.0530 $Y2=0.1510
r54 20 33 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1250 $X2=1.0530 $Y2=0.1400
r55 1 30 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=1.0530
+ $Y=0.1400 $X2=1.0530 $Y2=0.1400
r56 1 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.0530 $Y=0.1400
+ $X2=1.0530 $Y2=0.1400
r57 11 30 0.314665 $w=2.27e-07 $l=5e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.0530 $Y=0.1350 $X2=1.0530 $Y2=0.1400
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%SE VSS 34 5 6 8 13 7 11 9 12 2 1 10
c1 1 VSS 0.00182346f
c2 2 VSS 0.00390229f
c3 5 VSS 0.0426509f
c4 6 VSS 0.0814608f
c5 7 VSS 0.00156232f
c6 8 VSS 0.00027217f
c7 9 VSS 0.00480818f
c8 10 VSS 0.00504496f
c9 11 VSS 0.000202905f
c10 12 VSS 0.00563129f
c11 13 VSS 0.049185f
r1 1 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
r2 5 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r3 38 39 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2745
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r4 37 38 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2595
+ $Y=0.1350 $X2=0.2745 $Y2=0.1350
r5 36 37 0.699569 $w=1.3e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.1350 $X2=0.2595 $Y2=0.1350
r6 34 8 2.49951 $w=7.46154e-09 $l=1.95256e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.1340 $X2=0.2445 $Y2=0.1350
r7 8 36 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2445
+ $Y=0.1350 $X2=0.2565 $Y2=0.1350
r8 34 11 0.433689 $w=1.8e-08 $l=4.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.1340 $X2=0.2250 $Y2=0.1297
r9 11 32 3.53073 $w=1.4087e-08 $l=1.72e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.1297 $X2=0.2250 $Y2=0.1125
r10 10 28 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.2250 $Y=0.0360 $X2=0.2250
+ $Y2=0.0450
r11 31 32 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0900 $X2=0.2250 $Y2=0.1125
r12 30 31 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0675 $X2=0.2250 $Y2=0.0900
r13 7 30 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0495 $X2=0.2250 $Y2=0.0675
r14 7 28 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.2250 $Y=0.0495 $X2=0.2250
+ $Y2=0.0450
r15 7 10 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.0495 $X2=0.2250 $Y2=0.0360
r16 28 29 14.108 $w=1.3e-08 $l=6.05e-08 $layer=M2 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0450 $X2=0.2855 $Y2=0.0450
r17 26 29 109.716 $w=1.3e-08 $l=4.705e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.7560 $Y=0.0450 $X2=0.2855 $Y2=0.0450
r18 13 24 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=1.1905
+ $Y=0.0450 $X2=1.2150 $Y2=0.0450
r19 13 26 101.321 $w=1.3e-08 $l=4.345e-07 $layer=M2 $thickness=3.6e-08
+ $X=1.1905 $Y=0.0450 $X2=0.7560 $Y2=0.0450
r20 12 24 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=1.2150 $Y=0.0360 $X2=1.2150
+ $Y2=0.0450
r21 20 21 6.41272 $w=1.3e-08 $l=2.75e-08 $layer=M1 $thickness=3.6e-08 $X=1.2150
+ $Y=0.1085 $X2=1.2150 $Y2=0.1360
r22 19 20 8.51143 $w=1.3e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=1.2150
+ $Y=0.0720 $X2=1.2150 $Y2=0.1085
r23 9 19 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.2150
+ $Y=0.0495 $X2=1.2150 $Y2=0.0720
r24 9 12 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.2150 $Y=0.0495 $X2=1.2150 $Y2=0.0360
r25 9 24 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=1.2150 $Y=0.0495 $X2=1.2150
+ $Y2=0.0450
r26 6 2 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=1.2150
+ $Y=0.1350 $X2=1.2150 $Y2=0.1360
r27 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.2150 $Y=0.1360
+ $X2=1.2150 $Y2=0.1360
.ends

.subckt PM_SDFHx2_ASAP7_75t_R%CLKN VSS 13 14 15 72 74 26 7 22 17 16 19 21 1 8
+ 20 18 29 23 24 3 2 28 25 27
c1 1 VSS 0.00148421f
c2 2 VSS 0.000108839f
c3 3 VSS 0.000191685f
c4 7 VSS 0.00770043f
c5 8 VSS 0.0079155f
c6 13 VSS 0.0592771f
c7 14 VSS 0.0044842f
c8 15 VSS 0.00460295f
c9 16 VSS 0.00627171f
c10 17 VSS 0.00615507f
c11 18 VSS 0.0055848f
c12 19 VSS 0.00373678f
c13 20 VSS 0.00512251f
c14 21 VSS 0.00463376f
c15 22 VSS 0.000612442f
c16 23 VSS 0.000113531f
c17 24 VSS 0.000475371f
c18 25 VSS 0.00357059f
c19 26 VSS 0.00168129f
c20 27 VSS 0.00366918f
c21 28 VSS 0.00015415f
c22 29 VSS 0.0239372f
r1 74 73 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r2 17 73 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r3 72 71 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r4 16 71 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r5 8 69 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0550 $Y2=0.2340
r6 7 66 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0550 $Y2=0.0360
r7 68 69 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.2340 $X2=0.0550 $Y2=0.2340
r8 21 68 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0460 $Y2=0.2340
r9 21 27 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0180 $Y2=0.2340
r10 65 66 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.0360 $X2=0.0550 $Y2=0.0360
r11 20 65 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0460 $Y2=0.0360
r12 20 25 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0180 $Y2=0.0360
r13 27 62 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.2340 $X2=0.0180 $Y2=0.2125
r14 25 61 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.0360 $X2=0.0180 $Y2=0.0630
r15 1 56 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1440
r16 13 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r17 19 26 5.19594 $w=1.44151e-08 $l=2.80401e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1810 $X2=0.0165 $Y2=0.1530
r18 19 62 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1810 $X2=0.0180 $Y2=0.2125
r19 60 61 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0900 $X2=0.0180 $Y2=0.0630
r20 18 26 6.0121 $w=1.425e-08 $l=3.15357e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1215 $X2=0.0165 $Y2=0.1530
r21 18 60 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1215 $X2=0.0180 $Y2=0.0900
r22 2 50 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6210 $Y=0.1350
+ $X2=0.6210 $Y2=0.1395
r23 14 2 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1350
r24 22 56 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1235 $X2=0.1350 $Y2=0.1440
r25 53 54 1.90199 $w=1.38333e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.0255 $Y=0.1530 $X2=0.0345 $Y2=0.1530
r26 26 53 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0165
+ $Y=0.1530 $X2=0.0255 $Y2=0.1530
r27 28 50 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1620 $X2=0.6210 $Y2=0.1395
r28 28 41 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.6210 $Y=0.1620 $X2=0.6210
+ $Y2=0.1530
r29 23 50 5.47996 $w=1.3e-08 $l=2.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1160 $X2=0.6210 $Y2=0.1395
r30 48 49 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1530 $X2=0.1595 $Y2=0.1530
r31 48 56 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1350 $Y=0.1530
+ $X2=0.1350 $Y2=0.1440
r32 47 48 11.8927 $w=1.3e-08 $l=5.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.0840
+ $Y=0.1530 $X2=0.1350 $Y2=0.1530
r33 46 47 11.8927 $w=1.3e-08 $l=5.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.0330
+ $Y=0.1530 $X2=0.0840 $Y2=0.1530
r34 46 54 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.0330 $Y=0.1530
+ $X2=0.0345 $Y2=0.1530
r35 44 49 7.81186 $w=1.3e-08 $l=3.35e-08 $layer=M2 $thickness=3.6e-08 $X=0.1930
+ $Y=0.1530 $X2=0.1595 $Y2=0.1530
r36 43 44 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.2740
+ $Y=0.1530 $X2=0.1930 $Y2=0.1530
r37 41 42 15.2739 $w=1.3e-08 $l=6.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1530 $X2=0.6865 $Y2=0.1530
r38 41 50 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.6210 $Y=0.1530 $X2=0.6210
+ $Y2=0.1395
r39 40 41 34.1623 $w=1.3e-08 $l=1.465e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.4745 $Y=0.1530 $X2=0.6210 $Y2=0.1530
r40 40 43 46.7545 $w=1.3e-08 $l=2.005e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.4745 $Y=0.1530 $X2=0.2740 $Y2=0.1530
r41 29 39 18.3054 $w=1.3e-08 $l=7.85e-08 $layer=M2 $thickness=3.6e-08 $X=0.8125
+ $Y=0.1530 $X2=0.8910 $Y2=0.1530
r42 29 42 29.3819 $w=1.3e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.8125
+ $Y=0.1530 $X2=0.6865 $Y2=0.1530
r43 37 39 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.8910 $Y=0.1440
+ $X2=0.8910 $Y2=0.1530
r44 24 37 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1135 $X2=0.8910 $Y2=0.1440
r45 15 3 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.8910
+ $Y=0.1350 $X2=0.8910 $Y2=0.1350
r46 3 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8910 $Y=0.1350
+ $X2=0.8910 $Y2=0.1440
r47 8 17 1e-05
r48 7 16 1e-05
.ends


*
.SUBCKT SDFHx2_ASAP7_75t_R VSS VDD CLK SE D SI QN
*
* VSS VSS
* VDD VDD
* CLK CLK
* SE SE
* D D
* SI SI
* QN QN
*
*

MM20 N_MM20_d N_MM20_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM23 N_MM23_d N_MM22_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM0 N_MM0_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM28 N_MM28_d N_MM2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM29 N_MM29_d N_MM26_g N_MM29_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM27_g N_MM5_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM10_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM6 N_MM6_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM12 N_MM12_d N_MM12_g N_MM12_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM17 N_MM17_d N_MM17_g N_MM17_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM16 N_MM16_d N_MM16_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM14 N_MM14_d N_MM14_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM30 N_MM30_d N_MM30_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM24 N_MM24_d N_MM24_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@2 N_MM24@2_d N_MM24@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM21 N_MM21_d N_MM20_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM22 N_MM22_d N_MM22_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g N_MM3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM26 N_MM26_d N_MM26_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM27 N_MM27_d N_MM27_g N_MM27_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM13 N_MM13_d N_MM17_g N_MM13_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM18 N_MM18_d N_MM18_g N_MM18_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM19 N_MM19_d N_MM16_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM15 N_MM15_d N_MM14_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM31 N_MM31_d N_MM30_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM25 N_MM25_d N_MM24_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@2 N_MM25@2_d N_MM24@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "SDFHx2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "SDFHx2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_SDFHx2_ASAP7_75t_R%NET0167 VSS N_MM28_d N_MM29_s N_NET0167_1
+ PM_SDFHx2_ASAP7_75t_R%NET0167
cc_1 N_NET0167_1 N_MM2_g 0.0173478f
cc_2 N_NET0167_1 N_MM26_g 0.0172429f
x_PM_SDFHx2_ASAP7_75t_R%D VSS D N_MM26_g N_D_1 N_D_5 PM_SDFHx2_ASAP7_75t_R%D
cc_3 N_MM26_g N_SEN_16 0.000472394f
cc_4 N_MM26_g N_SEN_1 0.000865616f
cc_5 N_D_1 N_SEN_1 0.00120732f
cc_6 N_D_5 N_SEN_14 0.0015929f
cc_7 N_D N_SEN_12 0.00215936f
cc_8 N_MM26_g N_MM2_g 0.00504614f
x_PM_SDFHx2_ASAP7_75t_R%NET0166 VSS N_MM0_d N_MM5_s N_NET0166_7 N_NET0166_9
+ N_NET0166_1 N_NET0166_11 N_NET0166_12 N_NET0166_10 N_NET0166_8 N_NET0166_2
+ PM_SDFHx2_ASAP7_75t_R%NET0166
cc_9 N_NET0166_7 N_SE_1 0.00125798f
cc_10 N_NET0166_9 N_SE_10 0.000664406f
cc_11 N_NET0166_1 N_SE_8 0.0008353f
cc_12 N_NET0166_11 N_SE_7 0.00129003f
cc_13 N_NET0166_12 N_SE_10 0.00133749f
cc_14 N_NET0166_1 N_MM3_g 0.00158735f
cc_15 N_NET0166_11 N_SE_8 0.00366273f
cc_16 N_NET0166_10 N_SE_13 0.00425215f
cc_17 N_NET0166_7 N_MM3_g 0.0341298f
cc_18 N_NET0166_10 N_SEN_12 0.000325061f
cc_19 N_NET0166_10 N_SEN_16 0.000377331f
cc_20 N_NET0166_11 N_SEN_12 0.00111086f
cc_21 N_NET0166_10 N_SEN_14 0.00546734f
cc_22 N_NET0166_8 N_SI_1 0.00129825f
cc_23 N_NET0166_2 N_MM27_g 0.001532f
cc_24 N_NET0166_8 N_MM27_g 0.0348469f
x_PM_SDFHx2_ASAP7_75t_R%noxref_33 VSS N_noxref_33_1
+ PM_SDFHx2_ASAP7_75t_R%noxref_33
cc_25 N_noxref_33_1 N_MM30_g 0.00557958f
cc_26 N_noxref_33_1 N_SEN_3 0.00139286f
cc_27 N_noxref_33_1 N_SEN_10 0.0170312f
cc_28 N_noxref_33_1 N_SS_10 0.000446651f
cc_29 N_noxref_33_1 N_noxref_31_1 0.00768977f
cc_30 N_noxref_33_1 N_noxref_32_1 0.000507335f
x_PM_SDFHx2_ASAP7_75t_R%noxref_34 VSS N_noxref_34_1
+ PM_SDFHx2_ASAP7_75t_R%noxref_34
cc_31 N_noxref_34_1 N_MM30_g 0.00567945f
cc_32 N_noxref_34_1 N_SEN_4 0.000300671f
cc_33 N_noxref_34_1 N_SEN_11 0.0166867f
cc_34 N_noxref_34_1 N_SS_11 0.000611822f
cc_35 N_noxref_34_1 N_noxref_31_1 0.000510556f
cc_36 N_noxref_34_1 N_noxref_32_1 0.00786738f
cc_37 N_noxref_34_1 N_noxref_33_1 0.00152218f
x_PM_SDFHx2_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_SDFHx2_ASAP7_75t_R%noxref_24
cc_38 N_noxref_24_1 N_MM20_g 0.00369504f
cc_39 N_noxref_24_1 N_CLKN_26 5.78412e-20
cc_40 N_noxref_24_1 N_CLKN_25 5.79853e-20
cc_41 N_noxref_24_1 N_CLKN_19 6.56208e-20
cc_42 N_noxref_24_1 N_CLKN_18 0.000314669f
cc_43 N_noxref_24_1 N_CLKN_7 0.000504732f
cc_44 N_noxref_24_1 N_CLKN_16 0.0276257f
x_PM_SDFHx2_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_SDFHx2_ASAP7_75t_R%noxref_25
cc_45 N_noxref_25_1 N_MM20_g 0.00368577f
cc_46 N_noxref_25_1 N_CLKN_27 6.01554e-20
cc_47 N_noxref_25_1 N_CLKN_26 8.78806e-20
cc_48 N_noxref_25_1 N_CLKN_18 0.000151904f
cc_49 N_noxref_25_1 N_CLKN_19 0.000202276f
cc_50 N_noxref_25_1 N_CLKN_8 0.000500585f
cc_51 N_noxref_25_1 N_CLKN_17 0.0276135f
cc_52 N_noxref_25_1 N_noxref_24_1 0.00204371f
x_PM_SDFHx2_ASAP7_75t_R%PD4 VSS N_MM18_s N_MM19_d N_PD4_1
+ PM_SDFHx2_ASAP7_75t_R%PD4
cc_53 N_PD4_1 N_MM18_g 0.00783222f
cc_54 N_PD4_1 N_MM16_g 0.00773636f
x_PM_SDFHx2_ASAP7_75t_R%PD3 VSS N_MM9_s N_MM8_d N_PD3_1
+ PM_SDFHx2_ASAP7_75t_R%PD3
cc_55 N_PD3_1 N_MM9_g 0.00777478f
cc_56 N_PD3_1 N_MM11_g 0.0078334f
x_PM_SDFHx2_ASAP7_75t_R%CLK VSS CLK N_MM20_g N_CLK_4 N_CLK_6 N_CLK_1 N_CLK_5
+ PM_SDFHx2_ASAP7_75t_R%CLK
x_PM_SDFHx2_ASAP7_75t_R%SI VSS SI N_MM27_g N_SI_5 N_SI_1 N_SI_4 N_SI_6 N_SI_7
+ PM_SDFHx2_ASAP7_75t_R%SI
cc_57 N_SI_5 N_CLKN_29 0.00248803f
cc_58 N_SI_1 N_MM26_g 0.000900113f
cc_59 N_SI_4 N_D_5 0.00100829f
cc_60 N_MM27_g N_MM26_g 0.00404443f
x_PM_SDFHx2_ASAP7_75t_R%noxref_26 VSS N_noxref_26_1
+ PM_SDFHx2_ASAP7_75t_R%noxref_26
cc_61 N_noxref_26_1 N_MM22_g 0.00351361f
cc_62 N_noxref_26_1 N_CLKB_20 0.000144085f
cc_63 N_noxref_26_1 N_CLKB_6 0.00043246f
cc_64 N_noxref_26_1 N_CLKB_18 0.0270419f
cc_65 N_noxref_26_1 N_NET0166_7 0.000552006f
x_PM_SDFHx2_ASAP7_75t_R%noxref_28 VSS N_noxref_28_1
+ PM_SDFHx2_ASAP7_75t_R%noxref_28
cc_66 N_noxref_28_1 N_MM3_g 0.00161736f
cc_67 N_noxref_28_1 N_CLKB_6 9.95779e-20
cc_68 N_noxref_28_1 N_CLKB_18 0.0005185f
cc_69 N_noxref_28_1 N_NET0166_7 0.0359661f
cc_70 N_noxref_28_1 N_noxref_26_1 0.00769511f
cc_71 N_noxref_28_1 N_noxref_27_1 0.000469731f
x_PM_SDFHx2_ASAP7_75t_R%noxref_29 VSS N_noxref_29_1
+ PM_SDFHx2_ASAP7_75t_R%noxref_29
cc_72 N_noxref_29_1 N_MM3_g 0.00146625f
cc_73 N_noxref_29_1 N_CLKB_20 0.000107429f
cc_74 N_noxref_29_1 N_CLKB_19 0.000577319f
cc_75 N_noxref_29_1 N_NET0120_8 0.0360183f
cc_76 N_noxref_29_1 N_noxref_26_1 0.00046653f
cc_77 N_noxref_29_1 N_noxref_27_1 0.00771771f
cc_78 N_noxref_29_1 N_noxref_28_1 0.00123961f
x_PM_SDFHx2_ASAP7_75t_R%noxref_30 VSS N_noxref_30_1
+ PM_SDFHx2_ASAP7_75t_R%noxref_30
cc_79 N_noxref_30_1 N_MM27_g 0.00149574f
cc_80 N_noxref_30_1 N_SI_1 0.00244779f
cc_81 N_noxref_30_1 N_CLKB_1 0.000184852f
cc_82 N_noxref_30_1 N_MM1_g 0.010795f
cc_83 N_noxref_30_1 N_NET0120_2 0.00115771f
cc_84 N_noxref_30_1 N_NET0120_10 0.0161653f
cc_85 N_noxref_30_1 N_NET0120_9 0.0552353f
cc_86 N_noxref_30_1 N_NET0166_8 0.0370743f
x_PM_SDFHx2_ASAP7_75t_R%PD2 VSS N_MM10_s N_MM11_d N_PD2_4 N_PD2_5 N_PD2_1
+ PM_SDFHx2_ASAP7_75t_R%PD2
cc_87 N_PD2_4 N_MM10_g 0.0150098f
cc_88 N_PD2_4 N_CLKB_8 0.000126164f
cc_89 N_PD2_4 N_CLKB_2 0.000277591f
cc_90 N_PD2_5 N_CLKB_8 0.00167265f
cc_91 N_PD2_1 N_MM9_g 0.00209568f
cc_92 N_PD2_5 N_MM9_g 0.00734713f
cc_93 N_PD2_4 N_MM9_g 0.023831f
cc_94 N_PD2_5 N_MM11_g 0.0148551f
cc_95 N_PD2_4 N_MH_14 0.000321626f
cc_96 N_PD2_4 N_MH_3 0.000612784f
cc_97 N_PD2_1 N_MH_14 0.00347559f
x_PM_SDFHx2_ASAP7_75t_R%MH VSS N_MM7_g N_MM4_d N_MM9_d N_MM1_d N_MM10_d N_MH_10
+ N_MH_20 N_MH_14 N_MH_12 N_MH_16 N_MH_3 N_MH_4 N_MH_18 N_MH_17 N_MH_21 N_MH_1
+ N_MH_19 N_MH_15 PM_SDFHx2_ASAP7_75t_R%MH
cc_98 N_MH_10 N_CLKN_23 0.000252149f
cc_99 N_MH_10 N_CLKN_3 0.000109831f
cc_100 N_MH_10 N_MM17_g 0.000137083f
cc_101 N_MH_10 N_CLKN_28 0.000294078f
cc_102 N_MH_20 N_CLKN_28 0.000318978f
cc_103 N_MH_14 N_CLKN_28 0.000449092f
cc_104 N_MH_12 N_MM10_g 0.0163783f
cc_105 N_MH_16 N_CLKN_23 0.00052741f
cc_106 N_MH_3 N_CLKN_2 0.000605382f
cc_107 N_MH_4 N_CLKN_23 0.000808611f
cc_108 N_MH_18 N_CLKN_29 0.000903248f
cc_109 N_MH_4 N_MM10_g 0.00111183f
cc_110 N_MH_3 N_MM10_g 0.00122537f
cc_111 N_MH_10 N_CLKN_2 0.00160934f
cc_112 N_MH_17 N_CLKN_29 0.00166276f
cc_113 N_MH_17 N_CLKN_28 0.00211064f
cc_114 N_MH_10 N_MM10_g 0.0527294f
cc_115 N_MH_10 N_CLKB_21 0.00012272f
cc_116 N_MH_10 N_CLKB_22 0.00034123f
cc_117 N_MH_10 N_MM1_g 0.000428565f
cc_118 N_MH_10 N_CLKB_1 0.000203139f
cc_119 N_MH_3 N_CLKB_21 0.000340598f
cc_120 N_MH_3 N_CLKB_25 0.00035961f
cc_121 N_MH_21 N_CLKB_22 0.000404273f
cc_122 N_MH_17 N_CLKB_22 0.00646269f
cc_123 N_MH_17 N_CLKB_2 0.000497725f
cc_124 N_MH_1 N_CLKB_8 0.00208662f
cc_125 N_MH_4 N_MM9_g 0.000634f
cc_126 N_MH_12 N_CLKB_1 0.000668058f
cc_127 N_MH_17 N_CLKB_8 0.000774309f
cc_128 N_MH_14 N_CLKB_26 0.00141722f
cc_129 N_MH_18 N_CLKB_22 0.00150075f
cc_130 N_MH_3 N_MM1_g 0.00156427f
cc_131 N_MH_14 N_CLKB_25 0.00377685f
cc_132 N_MM7_g N_CLKB_8 0.00508852f
cc_133 N_MH_12 N_MM1_g 0.0330036f
cc_134 N_MM7_g N_MM12_g 0.0127442f
cc_135 N_MH_10 N_MM9_g 0.0361859f
cc_136 N_MH_19 N_MS_18 0.000267399f
cc_137 N_MH_4 N_MS_1 0.000360593f
cc_138 N_MH_18 N_MS_19 0.000374126f
cc_139 N_MH_18 N_MS_1 0.000663171f
cc_140 N_MM7_g N_MS_3 0.000938193f
cc_141 N_MH_18 N_MS_17 0.000995644f
cc_142 N_MH_1 N_MS_14 0.0010038f
cc_143 N_MH_1 N_MS_1 0.00130311f
cc_144 N_MM7_g N_MS_12 0.00632838f
cc_145 N_MM7_g N_MS_1 0.00241402f
cc_146 N_MM7_g N_MS_11 0.00639821f
cc_147 N_MH_18 N_MS_14 0.00459509f
cc_148 N_MH_16 N_MS_18 0.00497709f
cc_149 N_MM7_g N_MM11_g 0.0294176f
x_PM_SDFHx2_ASAP7_75t_R%noxref_27 VSS N_noxref_27_1
+ PM_SDFHx2_ASAP7_75t_R%noxref_27
cc_150 N_noxref_27_1 N_MM22_g 0.00353333f
cc_151 N_noxref_27_1 N_CLKB_20 0.000174169f
cc_152 N_noxref_27_1 N_CLKB_7 0.000434949f
cc_153 N_noxref_27_1 N_CLKB_19 0.026989f
cc_154 N_noxref_27_1 N_NET0120_8 0.000588846f
cc_155 N_noxref_27_1 N_noxref_26_1 0.00148613f
x_PM_SDFHx2_ASAP7_75t_R%NET0141 VSS N_MM3_s N_MM2_d N_MM26_d N_MM27_s
+ N_NET0141_7 N_NET0141_9 N_NET0141_1 N_NET0141_2 N_NET0141_8
+ PM_SDFHx2_ASAP7_75t_R%NET0141
cc_156 N_NET0141_7 N_SE_1 0.000978466f
cc_157 N_NET0141_9 N_SE_8 0.0006848f
cc_158 N_NET0141_1 N_MM3_g 0.000836137f
cc_159 N_NET0141_7 N_MM3_g 0.0329628f
cc_160 N_NET0141_7 N_SEN_1 0.000921232f
cc_161 N_NET0141_1 N_MM2_g 0.000852895f
cc_162 N_NET0141_9 N_SEN_12 0.00218874f
cc_163 N_NET0141_7 N_MM2_g 0.033024f
cc_164 N_NET0141_2 N_MM26_g 0.000866208f
cc_165 N_NET0141_9 N_D 0.00225353f
cc_166 N_NET0141_8 N_MM26_g 0.0340439f
cc_167 N_NET0141_9 N_SI_4 0.000662024f
cc_168 N_NET0141_8 N_SI_1 0.000778003f
cc_169 N_NET0141_2 N_MM27_g 0.000816974f
cc_170 N_NET0141_8 N_MM27_g 0.0335805f
cc_171 N_NET0141_9 N_CLKB_26 0.00296816f
cc_172 N_NET0141_2 N_NET0120_11 0.000548151f
cc_173 N_NET0141_7 N_NET0120_8 0.00110581f
cc_174 N_NET0141_8 N_NET0120_9 0.000555219f
cc_175 N_NET0141_1 N_NET0120_11 0.000597971f
cc_176 N_NET0141_8 N_NET0120_2 0.00130088f
cc_177 N_NET0141_2 N_NET0120_2 0.00161278f
cc_178 N_NET0141_1 N_NET0120_1 0.00303227f
cc_179 N_NET0141_9 N_NET0120_11 0.0131795f
x_PM_SDFHx2_ASAP7_75t_R%MS VSS N_MM11_g N_MM6_d N_MM12_d N_MM7_d N_MM13_d
+ N_MS_13 N_MS_17 N_MS_19 N_MS_18 N_MS_3 N_MS_15 N_MS_12 N_MS_1 N_MS_11 N_MS_4
+ N_MS_14 N_MS_16 PM_SDFHx2_ASAP7_75t_R%MS
cc_180 N_MS_13 N_CLKN_24 0.000245511f
cc_181 N_MS_13 N_MM10_g 0.000137844f
cc_182 N_MS_13 N_CLKN_29 0.000349468f
cc_183 N_MS_13 N_CLKN_3 0.000222252f
cc_184 N_MS_17 N_CLKN_24 0.0045445f
cc_185 N_MS_17 N_CLKN_3 0.000289706f
cc_186 N_MS_19 N_CLKN_24 0.000418989f
cc_187 N_MS_18 N_CLKN_29 0.00162458f
cc_188 N_MS_13 N_MM17_g 0.0155046f
cc_189 N_MS_18 N_SEN_16 0.000925052f
cc_190 N_MS_19 N_SEN_16 0.00303695f
cc_191 N_MS_3 N_CLKB_22 0.00014273f
cc_192 N_MS_3 N_CLKB_8 0.000652432f
cc_193 N_MS_3 N_CLKB_2 9.25654e-20
cc_194 N_MS_3 N_CLKB_26 0.000142224f
cc_195 N_MS_15 N_CLKB_22 0.000281055f
cc_196 N_MS_13 N_MM12_g 0.00786932f
cc_197 N_MS_15 N_CLKB_8 0.000361999f
cc_198 N_MS_12 N_MM12_g 0.00781547f
cc_199 N_MS_1 N_MM9_g 0.000704144f
cc_200 N_MS_17 N_CLKB_8 0.00154178f
cc_201 N_MS_11 N_MM12_g 0.006509f
cc_202 N_MS_4 N_MM12_g 0.00257216f
cc_203 N_MS_4 N_CLKB_8 0.00639183f
cc_204 N_MM11_g N_MM9_g 0.0141679f
cc_205 N_MS_3 N_MM12_g 0.0259814f
x_PM_SDFHx2_ASAP7_75t_R%NET0120 VSS N_MM3_d N_MM27_d N_MM1_s N_NET0120_8
+ N_NET0120_1 N_NET0120_2 N_NET0120_9 N_NET0120_11 N_NET0120_10
+ PM_SDFHx2_ASAP7_75t_R%NET0120
cc_206 N_NET0120_8 N_SE_8 0.000715972f
cc_207 N_NET0120_8 N_SE_1 0.00100337f
cc_208 N_NET0120_1 N_MM3_g 0.0013145f
cc_209 N_NET0120_8 N_MM3_g 0.0341033f
cc_210 N_NET0120_2 N_SI_5 0.00063876f
cc_211 N_NET0120_9 N_SI_1 0.00143546f
cc_212 N_NET0120_2 N_SI_6 0.00293469f
cc_213 N_NET0120_11 N_SI_6 0.00312868f
cc_214 N_NET0120_9 N_MM27_g 0.0350051f
cc_215 N_NET0120_10 N_CLKB_20 4.87542e-20
cc_216 N_NET0120_10 N_CLKB_24 0.00028648f
cc_217 N_NET0120_10 N_CLKB_7 0.000132986f
cc_218 N_NET0120_10 N_CLKB_19 0.000143194f
cc_219 N_NET0120_10 N_CLKB_1 0.00101257f
cc_220 N_NET0120_10 N_CLKB_25 0.000340289f
cc_221 N_NET0120_10 N_CLKB_21 0.000351433f
cc_222 N_NET0120_1 N_CLKB_20 0.000922357f
cc_223 N_NET0120_2 N_MM1_g 0.00158943f
cc_224 N_NET0120_11 N_CLKB_26 0.00368542f
cc_225 N_NET0120_10 N_MM1_g 0.0338943f
cc_226 N_NET0120_2 N_MH_3 0.00118827f
cc_227 N_NET0120_2 N_MH_12 0.00290416f
x_PM_SDFHx2_ASAP7_75t_R%NET0118 VSS N_MM29_d N_MM5_d N_MM4_s N_NET0118_8
+ N_NET0118_9 N_NET0118_2 N_NET0118_7 N_NET0118_1 PM_SDFHx2_ASAP7_75t_R%NET0118
cc_228 N_NET0118_8 N_CLKN_2 0.000897591f
cc_229 N_NET0118_9 N_CLKN_23 0.000742631f
cc_230 N_NET0118_2 N_MM10_g 0.000866236f
cc_231 N_NET0118_9 N_CLKN_29 0.000921737f
cc_232 N_NET0118_8 N_MM10_g 0.0327391f
cc_233 N_NET0118_9 N_SE_13 0.00227238f
cc_234 N_NET0118_9 N_MM2_g 0.000310008f
cc_235 N_NET0118_9 N_SEN_12 0.000111392f
cc_236 N_NET0118_9 N_SEN_14 0.000544193f
cc_237 N_NET0118_9 N_SEN_16 0.00391671f
cc_238 N_NET0118_7 N_D_1 0.000880932f
cc_239 N_NET0118_1 N_MM26_g 0.00126279f
cc_240 N_NET0118_9 N_D_5 0.00271958f
cc_241 N_NET0118_7 N_MM26_g 0.0342531f
cc_242 N_NET0118_9 N_SI_4 0.000432257f
cc_243 N_NET0118_1 N_MM27_g 0.000757283f
cc_244 N_NET0118_7 N_SI_1 0.000820405f
cc_245 N_NET0118_9 N_SI_7 0.00250569f
cc_246 N_NET0118_7 N_MM27_g 0.033464f
cc_247 N_NET0118_8 N_CLKB_21 0.000153127f
cc_248 N_NET0118_8 N_CLKB_1 0.00111444f
cc_249 N_NET0118_2 N_MM1_g 0.00116662f
cc_250 N_NET0118_9 N_CLKB_21 0.00236428f
cc_251 N_NET0118_8 N_MM1_g 0.0355577f
cc_252 N_NET0118_8 N_MH_10 0.00114786f
cc_253 N_NET0118_9 N_MH_15 0.000948568f
cc_254 N_NET0118_2 N_MH_4 0.0036769f
cc_255 N_NET0118_7 N_NET0166_10 0.000583281f
cc_256 N_NET0118_9 N_NET0166_2 0.000634274f
cc_257 N_NET0118_7 N_NET0166_8 0.000642339f
cc_258 N_NET0118_1 N_NET0166_2 0.00381284f
cc_259 N_NET0118_9 N_NET0166_10 0.00907244f
x_PM_SDFHx2_ASAP7_75t_R%noxref_31 VSS N_noxref_31_1
+ PM_SDFHx2_ASAP7_75t_R%noxref_31
cc_260 N_noxref_31_1 N_SEN_3 0.00116295f
cc_261 N_noxref_31_1 N_SS_10 0.0170021f
cc_262 N_noxref_31_1 N_MM14_g 0.0057463f
x_PM_SDFHx2_ASAP7_75t_R%SEN VSS N_MM2_g N_MM30_d N_MM31_d N_SEN_16 N_SEN_12
+ N_SEN_13 N_SEN_4 N_SEN_10 N_SEN_11 N_SEN_14 N_SEN_3 N_SEN_1 N_SEN_15
+ PM_SDFHx2_ASAP7_75t_R%SEN
cc_263 N_SEN_16 N_CLKN_24 0.00295696f
cc_264 N_SEN_16 N_CLKN_23 0.000503602f
cc_265 N_SEN_12 N_CLKN_29 0.00327767f
cc_266 N_SEN_16 N_CLKN_29 0.0107458f
cc_267 N_SEN_13 N_SE_9 0.00808565f
cc_268 N_SEN_4 N_SE_9 0.000213952f
cc_269 N_SEN_10 N_MM30_g 0.023221f
cc_270 N_SEN_11 N_MM30_g 0.00679819f
cc_271 N_SEN_14 N_SE_13 0.000247294f
cc_272 N_SEN_3 N_SE_9 0.000259952f
cc_273 N_SEN_1 N_SE_8 0.000309112f
cc_274 N_SEN_13 N_SE_12 0.000329572f
cc_275 N_SEN_4 N_MM30_g 0.00034942f
cc_276 N_SEN_3 N_SE_2 0.000410532f
cc_277 N_SEN_15 N_SE_9 0.000417746f
cc_278 N_SEN_13 N_SE_2 0.000422053f
cc_279 N_SEN_1 N_SE_1 0.00125681f
cc_280 N_SEN_12 N_SE_13 0.000479966f
cc_281 N_SEN_13 N_SE_13 0.000514992f
cc_282 N_SEN_3 N_MM30_g 0.00093838f
cc_283 N_SEN_12 N_SE_8 0.00172568f
cc_284 N_MM2_g N_MM3_g 0.00330887f
cc_285 N_SEN_16 N_SE_13 0.0644899f
x_PM_SDFHx2_ASAP7_75t_R%noxref_35 VSS N_noxref_35_1
+ PM_SDFHx2_ASAP7_75t_R%noxref_35
cc_286 N_noxref_35_1 N_MM24@2_g 0.00150406f
cc_287 N_noxref_35_1 N_QN_7 0.000832913f
x_PM_SDFHx2_ASAP7_75t_R%QN VSS QN N_MM24_d N_MM24@2_d N_MM25_d N_MM25@2_d
+ N_QN_9 N_QN_7 N_QN_8 N_QN_10 N_QN_11 N_QN_1 N_QN_2 PM_SDFHx2_ASAP7_75t_R%QN
cc_288 N_QN_9 N_SE_9 0.000631852f
cc_289 N_QN_9 N_SE_13 0.000267986f
cc_290 N_QN_9 N_SE_12 0.00158178f
cc_291 N_QN_7 N_SH_21 0.000914892f
cc_292 N_QN_7 N_SH_2 0.000443718f
cc_293 N_QN_7 N_SH_26 0.000626944f
cc_294 N_QN_8 N_MM24_g 0.0308852f
cc_295 N_QN_10 N_SH_21 0.000955777f
cc_296 N_QN_11 N_SH_2 0.00118399f
cc_297 N_QN_1 N_MM24_g 0.00205448f
cc_298 N_QN_2 N_SH_21 0.00241359f
cc_299 N_QN_2 N_MM24_g 0.00243743f
cc_300 N_QN_8 N_SH_2 0.00460238f
cc_301 N_QN_7 N_MM24@2_g 0.0372062f
cc_302 N_QN_7 N_MM24_g 0.0681535f
x_PM_SDFHx2_ASAP7_75t_R%noxref_36 VSS N_noxref_36_1
+ PM_SDFHx2_ASAP7_75t_R%noxref_36
cc_303 N_noxref_36_1 N_MM24@2_g 0.00150783f
cc_304 N_noxref_36_1 N_QN_8 0.000826366f
cc_305 N_noxref_36_1 N_noxref_35_1 0.00177706f
x_PM_SDFHx2_ASAP7_75t_R%PD5 VSS N_MM17_s N_MM16_d N_PD5_4 N_PD5_1 N_PD5_5
+ PM_SDFHx2_ASAP7_75t_R%PD5
cc_306 N_PD5_4 N_MM17_g 0.0152551f
cc_307 N_PD5_1 N_MM18_g 0.000757612f
cc_308 N_PD5_5 N_MM18_g 0.00693338f
cc_309 N_PD5_4 N_MM18_g 0.0239646f
cc_310 N_PD5_1 N_MM16_g 0.000892078f
cc_311 N_PD5_5 N_MM16_g 0.0155996f
cc_312 N_PD5_1 N_SH_14 0.000514885f
cc_313 N_PD5_1 N_SH_16 0.000490453f
cc_314 N_PD5_1 N_SH_17 0.000570902f
cc_315 N_PD5_4 N_SH_5 0.000658081f
cc_316 N_PD5_1 N_SH_23 0.00237847f
x_PM_SDFHx2_ASAP7_75t_R%noxref_32 VSS N_noxref_32_1
+ PM_SDFHx2_ASAP7_75t_R%noxref_32
cc_317 N_noxref_32_1 N_SEN_11 0.000618213f
cc_318 N_noxref_32_1 N_SS_11 0.0170395f
cc_319 N_noxref_32_1 N_MM14_g 0.00582072f
cc_320 N_noxref_32_1 N_noxref_31_1 0.00153605f
x_PM_SDFHx2_ASAP7_75t_R%CLKB VSS N_MM1_g N_MM9_g N_MM12_g N_MM18_g N_MM23_d
+ N_MM22_d N_CLKB_26 N_CLKB_19 N_CLKB_7 N_CLKB_18 N_CLKB_24 N_CLKB_6 N_CLKB_20
+ N_CLKB_23 N_CLKB_4 N_CLKB_22 N_CLKB_21 N_CLKB_8 N_CLKB_2 N_CLKB_1 N_CLKB_25
+ PM_SDFHx2_ASAP7_75t_R%CLKB
cc_321 N_CLKB_26 N_CLK_5 5.25347e-20
cc_322 N_CLKB_19 N_CLK_5 7.11297e-20
cc_323 N_CLKB_7 N_CLK_5 0.000491718f
cc_324 N_CLKB_18 N_CLK_5 8.91394e-20
cc_325 N_CLKB_24 N_CLK_5 0.000113024f
cc_326 N_CLKB_6 N_CLK_5 0.000386069f
cc_327 N_CLKB_20 N_CLK_6 0.000427282f
cc_328 N_CLKB_23 N_CLK_5 0.00187738f
cc_329 N_CLKB_23 N_CLKN_29 2.90609e-20
cc_330 N_CLKB_24 N_CLKN_29 3.70642e-20
cc_331 N_CLKB_23 N_CLKN_18 4.16972e-20
cc_332 N_CLKB_6 N_MM22_g 0.000651679f
cc_333 N_CLKB_24 N_CLKN_21 9.69708e-20
cc_334 N_CLKB_7 N_MM22_g 0.000788053f
cc_335 N_CLKB_4 N_MM17_g 0.000208159f
cc_336 N_CLKB_23 N_CLKN_22 0.000268624f
cc_337 N_CLKB_22 N_CLKN_29 0.000676953f
cc_338 N_CLKB_21 N_CLKN_29 0.00032759f
cc_339 N_CLKB_20 N_CLKN_22 0.00454098f
cc_340 N_CLKB_24 N_CLKN_22 0.000383004f
cc_341 N_CLKB_18 N_MM22_g 0.0386421f
cc_342 N_CLKB_19 N_MM22_g 0.0111504f
cc_343 N_CLKB_26 N_CLKN_23 0.000478614f
cc_344 N_CLKB_20 N_CLKN_29 0.00052875f
cc_345 N_CLKB_8 N_CLKN_24 0.000531969f
cc_346 N_CLKB_2 N_MM10_g 0.000560153f
cc_347 N_CLKB_20 N_CLKN_1 0.000579205f
cc_348 N_CLKB_8 N_CLKN_3 0.0027913f
cc_349 N_CLKB_19 N_CLKN_1 0.000784303f
cc_350 N_CLKB_1 N_CLKN_2 0.00222254f
cc_351 N_CLKB_25 N_CLKN_28 0.00165668f
cc_352 N_CLKB_21 N_CLKN_23 0.00265808f
cc_353 N_MM9_g N_MM10_g 0.00370403f
cc_354 N_CLKB_8 N_MM17_g 0.00493087f
cc_355 N_MM18_g N_MM17_g 0.00578287f
cc_356 N_MM1_g N_MM10_g 0.00704193f
cc_357 N_MM12_g N_MM17_g 0.0182753f
cc_358 N_CLKB_26 N_CLKN_29 0.0447356f
cc_359 N_CLKB_7 N_SE_11 4.71947e-20
cc_360 N_CLKB_6 N_SE_10 5.44479e-20
cc_361 N_MM18_g N_SE_13 0.000110728f
cc_362 N_CLKB_6 N_SE_7 0.000174715f
cc_363 N_CLKB_26 N_SE_13 0.000251283f
cc_364 N_CLKB_20 N_SE_7 0.00298567f
cc_365 N_CLKB_21 N_SE_13 0.000837113f
cc_366 N_CLKB_26 N_SE_8 0.00121828f
cc_367 N_CLKB_23 N_SE_10 0.00174526f
cc_368 N_CLKB_20 N_SE_11 0.00644922f
cc_369 N_MM1_g N_SI_5 7.57729e-20
cc_370 N_CLKB_1 N_SI_5 0.000390057f
cc_371 N_CLKB_26 N_SI_5 0.000985897f
cc_372 N_CLKB_26 N_SI_6 0.000321463f
cc_373 N_CLKB_21 N_SI_7 0.000812248f
cc_374 N_CLKB_25 N_SI_6 0.000920349f
cc_375 N_CLKB_21 N_SI_5 0.00266998f
x_PM_SDFHx2_ASAP7_75t_R%SS VSS N_MM16_g N_MM14_d N_MM15_d N_SS_14 N_SS_13
+ N_SS_12 N_SS_17 N_SS_16 N_SS_3 N_SS_4 N_SS_15 N_SS_1 N_SS_10 N_SS_11
+ PM_SDFHx2_ASAP7_75t_R%SS
cc_376 N_SS_14 N_SE_13 0.000528557f
cc_377 N_SS_13 N_SE_13 0.000906364f
cc_378 N_SS_12 N_SE_13 0.0029651f
cc_379 N_SS_14 N_SEN_3 0.00123036f
cc_380 N_SS_14 N_SEN_4 0.000106637f
cc_381 N_SS_14 N_SEN_15 0.000108856f
cc_382 N_SS_13 N_SEN_16 0.00035578f
cc_383 N_SS_17 N_SEN_13 0.000424246f
cc_384 N_SS_16 N_SEN_15 0.000788228f
cc_385 N_SS_12 N_SEN_16 0.00262149f
cc_386 N_SS_14 N_SEN_13 0.00845499f
cc_387 N_MM16_g N_CLKB_8 0.000681351f
cc_388 N_MM16_g N_CLKB_4 0.000426619f
cc_389 N_MM16_g N_MM18_g 0.0133591f
x_PM_SDFHx2_ASAP7_75t_R%SH VSS N_MM14_g N_MM24_g N_MM24@2_g N_MM13_s N_MM18_d
+ N_MM12_s N_MM17_d N_SH_6 N_SH_14 N_SH_15 N_SH_22 N_SH_16 N_SH_24 N_SH_18
+ N_SH_17 N_SH_5 N_SH_26 N_SH_21 N_SH_2 N_SH_23 N_SH_1 N_SH_19 N_SH_20 N_SH_25
+ PM_SDFHx2_ASAP7_75t_R%SH
cc_390 N_SH_6 N_MM17_g 0.000158318f
cc_391 N_SH_14 N_MM17_g 0.00676966f
cc_392 N_SH_15 N_MM17_g 0.00683991f
cc_393 N_SH_22 N_CLKN_24 0.000285603f
cc_394 N_SH_16 N_CLKN_24 0.000369687f
cc_395 N_SH_24 N_CLKN_24 0.000402567f
cc_396 N_SH_18 N_CLKN_24 0.000478144f
cc_397 N_SH_17 N_CLKN_3 0.000570191f
cc_398 N_SH_5 N_CLKN_3 0.000576027f
cc_399 N_SH_26 N_CLKN_29 0.000779023f
cc_400 N_SH_17 N_CLKN_24 0.00451947f
cc_401 N_SH_16 N_CLKN_29 0.00111364f
cc_402 N_SH_5 N_MM17_g 0.0183294f
cc_403 N_SH_21 N_SE_12 0.000229657f
cc_404 N_SH_17 N_SE_13 0.000315749f
cc_405 N_SH_2 N_SE_2 0.00162146f
cc_406 N_SH_16 N_SE_13 0.00102205f
cc_407 N_SH_26 N_SE_13 0.00209908f
cc_408 N_SH_23 N_SE_13 0.00268191f
cc_409 N_MM24_g N_MM30_g 0.00337225f
cc_410 N_SH_21 N_SE_9 0.00618393f
cc_411 N_SH_1 N_SEN_13 0.00014553f
cc_412 N_MM24_g N_SEN_3 7.12209e-20
cc_413 N_SH_19 N_SEN_16 0.000109197f
cc_414 N_SH_26 N_SEN_15 0.000118258f
cc_415 N_SH_21 N_SEN_13 0.000155127f
cc_416 N_SH_26 N_SEN_13 0.00158073f
cc_417 N_SH_21 N_SEN_15 0.000259176f
cc_418 N_SH_20 N_SEN_16 0.000283404f
cc_419 N_SH_16 N_SEN_16 0.000373784f
cc_420 N_SH_26 N_SEN_16 0.00458123f
cc_421 N_SH_17 N_SEN_16 0.00612084f
cc_422 N_SH_15 N_CLKB_8 8.1806e-20
cc_423 N_SH_15 N_CLKB_26 8.30648e-20
cc_424 N_MM14_g N_MM18_g 8.8363e-20
cc_425 N_SH_22 N_CLKB_8 0.000196954f
cc_426 N_SH_24 N_CLKB_8 0.000203975f
cc_427 N_SH_14 N_MM12_g 0.00680288f
cc_428 N_SH_6 N_CLKB_8 0.000276295f
cc_429 N_SH_19 N_CLKB_8 0.000396208f
cc_430 N_SH_17 N_CLKB_8 0.000448364f
cc_431 N_SH_18 N_CLKB_8 0.000562994f
cc_432 N_SH_15 N_CLKB_4 0.000673075f
cc_433 N_SH_6 N_MM18_g 0.00100239f
cc_434 N_SH_5 N_CLKB_8 0.00282998f
cc_435 N_SH_5 N_MM12_g 0.00947937f
cc_436 N_SH_15 N_MM18_g 0.0159993f
cc_437 N_SH_18 N_MS_3 9.84547e-20
cc_438 N_SH_22 N_MS_3 0.000179155f
cc_439 N_SH_15 N_MS_3 0.000436412f
cc_440 N_SH_6 N_MS_3 0.000220896f
cc_441 N_SH_14 N_MS_3 0.000232021f
cc_442 N_SH_14 N_MS_11 0.000234022f
cc_443 N_SH_22 N_MS_4 0.000335705f
cc_444 N_SH_6 N_MS_4 0.000424812f
cc_445 N_SH_16 N_MS_16 0.00043823f
cc_446 N_SH_22 N_MS_17 0.000517696f
cc_447 N_SH_15 N_MS_4 0.00059315f
cc_448 N_SH_16 N_MS_19 0.00132439f
cc_449 N_SH_5 N_MS_3 0.00373413f
cc_450 N_SH_18 N_MM16_g 0.000104039f
cc_451 N_SH_20 N_SS_13 0.000311072f
cc_452 N_MM14_g N_SS_3 0.000322891f
cc_453 N_MM14_g N_SS_4 0.00042065f
cc_454 N_SH_23 N_SS_15 0.000580125f
cc_455 N_SH_25 N_SS_16 0.000641443f
cc_456 N_SH_25 N_SS_14 0.00069774f
cc_457 N_SH_17 N_SS_1 0.000810777f
cc_458 N_SH_1 N_SS_14 0.000948913f
cc_459 N_MM14_g N_SS_1 0.00111318f
cc_460 N_SH_1 N_MM16_g 0.00135492f
cc_461 N_SH_19 N_SS_12 0.00154855f
cc_462 N_SH_26 N_SS_14 0.00169901f
cc_463 N_MM14_g N_SS_10 0.00649593f
cc_464 N_MM14_g N_SS_11 0.00660056f
cc_465 N_SH_17 N_SS_12 0.00462671f
cc_466 N_SH_20 N_SS_14 0.00484973f
cc_467 N_MM14_g N_MM16_g 0.0300221f
x_PM_SDFHx2_ASAP7_75t_R%SE VSS SE N_MM3_g N_MM30_g N_SE_8 N_SE_13 N_SE_7
+ N_SE_11 N_SE_9 N_SE_12 N_SE_2 N_SE_1 N_SE_10 PM_SDFHx2_ASAP7_75t_R%SE
cc_468 N_SE_8 N_CLKN_22 3.25212e-20
cc_469 N_SE_13 N_CLKN_23 3.39836e-20
cc_470 N_SE_7 N_CLKN_18 3.51134e-20
cc_471 N_SE_11 N_CLKN_1 3.66514e-20
cc_472 N_SE_11 N_CLKN_22 5.50724e-20
cc_473 N_SE_7 N_CLKN_29 0.000403674f
cc_474 N_SE_11 N_CLKN_29 0.000313663f
cc_475 N_SE_13 N_CLKN_24 0.000502662f
cc_476 N_SE_13 N_CLKN_29 0.00246309f
cc_477 N_SE_8 N_CLKN_29 0.00355184f
x_PM_SDFHx2_ASAP7_75t_R%CLKN VSS N_MM22_g N_MM10_g N_MM17_g N_MM20_d N_MM21_d
+ N_CLKN_26 N_CLKN_7 N_CLKN_22 N_CLKN_17 N_CLKN_16 N_CLKN_19 N_CLKN_21 N_CLKN_1
+ N_CLKN_8 N_CLKN_20 N_CLKN_18 N_CLKN_29 N_CLKN_23 N_CLKN_24 N_CLKN_3 N_CLKN_2
+ N_CLKN_28 N_CLKN_25 N_CLKN_27 PM_SDFHx2_ASAP7_75t_R%CLKN
cc_478 N_CLKN_26 N_MM20_g 0.000235536f
cc_479 N_CLKN_7 N_MM20_g 0.00109794f
cc_480 N_CLKN_22 N_MM20_g 0.000270134f
cc_481 N_CLKN_17 N_MM20_g 0.011216f
cc_482 N_CLKN_16 N_MM20_g 0.011219f
cc_483 N_CLKN_19 N_CLK_4 0.000475848f
cc_484 N_CLKN_21 N_CLK_4 0.000489228f
cc_485 N_CLKN_1 N_CLK_6 0.000644362f
cc_486 N_CLKN_8 N_MM20_g 0.000752868f
cc_487 N_CLKN_26 N_CLK_1 0.000930979f
cc_488 N_CLKN_20 N_CLK_6 0.000991634f
cc_489 N_CLKN_22 N_CLK_6 0.00104499f
cc_490 N_CLKN_18 N_CLK_6 0.00109856f
cc_491 N_CLKN_29 N_CLK_6 0.00130052f
cc_492 N_CLKN_22 N_CLK_4 0.00147124f
cc_493 N_CLKN_20 N_CLK_5 0.00188064f
cc_494 N_CLKN_1 N_CLK_1 0.002428f
cc_495 N_CLKN_26 N_CLK_4 0.00645141f
cc_496 N_MM22_g N_MM20_g 0.0351967f
*END of SDFHx2_ASAP7_75t_R.pxi
.ENDS
** Design:	SDFHx3_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "SDFHx3_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "SDFHx3_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_SDFHx3_ASAP7_75t_R%NET137 VSS 2 3 1
c1 1 VSS 0.000995612f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3780 $Y2=0.0675
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%noxref_33 VSS 1
c1 1 VSS 0.00365548f
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%noxref_34 VSS 1
c1 1 VSS 0.00399544f
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.00421237f
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.00426883f
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%noxref_31 VSS 1
c1 1 VSS 0.00360544f
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%noxref_32 VSS 1
c1 1 VSS 0.00379701f
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%NET134 VSS 14 27 7 9 1 11 12 10 8 2
c1 1 VSS 0.00638283f
c2 2 VSS 0.00557085f
c3 7 VSS 0.00466657f
c4 8 VSS 0.00320522f
c5 9 VSS 0.000876754f
c6 10 VSS 0.017526f
c7 11 VSS 0.00131496f
c8 12 VSS 0.00207232f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0675 $X2=0.4840 $Y2=0.0675
r2 27 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4715 $Y2=0.0675
r3 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0675
+ $X2=0.4860 $Y2=0.0360
r4 23 24 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4475
+ $Y=0.0360 $X2=0.4860 $Y2=0.0360
r5 22 23 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4070
+ $Y=0.0360 $X2=0.4475 $Y2=0.0360
r6 21 22 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.3875
+ $Y=0.0360 $X2=0.4070 $Y2=0.0360
r7 20 21 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3605
+ $Y=0.0360 $X2=0.3875 $Y2=0.0360
r8 19 20 7.92845 $w=1.3e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3265
+ $Y=0.0360 $X2=0.3605 $Y2=0.0360
r9 10 12 1.03257 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3085 $Y=0.0360 $X2=0.2970 $Y2=0.0360
r10 10 19 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3085
+ $Y=0.0360 $X2=0.3265 $Y2=0.0360
r11 12 18 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.2970 $Y2=0.0540
r12 9 17 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0720 $X2=0.2970 $Y2=0.0900
r13 9 18 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0720 $X2=0.2970 $Y2=0.0540
r14 16 17 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2835 $Y=0.0900 $X2=0.2970 $Y2=0.0900
r15 11 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0900 $X2=0.2835 $Y2=0.0900
r16 11 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0900
+ $X2=0.2700 $Y2=0.0945
r17 1 15 23.8708 $w=2.02e-08 $l=4.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.2700 $Y=0.0540 $X2=0.2700 $Y2=0.0945
r18 14 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r19 7 13 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r20 1 7 1e-05
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%noxref_35 VSS 1
c1 1 VSS 0.00540821f
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%noxref_36 VSS 1
c1 1 VSS 0.00534632f
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%QN VSS 32 24 25 35 42 43 45 13 19 3 15 4 18 1 2
+ 16 14
c1 1 VSS 0.0107234f
c2 2 VSS 0.0103551f
c3 3 VSS 0.00786439f
c4 4 VSS 0.00791459f
c5 13 VSS 0.0046069f
c6 14 VSS 0.00345509f
c7 15 VSS 0.00454213f
c8 16 VSS 0.00344276f
c9 17 VSS 0.0149105f
c10 18 VSS 0.0142565f
c11 19 VSS 0.00383404f
c12 20 VSS 0.00279963f
c13 21 VSS 0.00285696f
r1 16 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.3895 $Y=0.2025 $X2=1.4020 $Y2=0.2025
r2 45 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.3870 $Y=0.2025 $X2=1.3895 $Y2=0.2025
r3 43 41 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.3130 $Y=0.2025 $X2=1.3105 $Y2=0.2025
r4 2 41 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.2960 $Y=0.2025 $X2=1.3105 $Y2=0.2025
r5 15 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.2815 $Y=0.2025 $X2=1.2960 $Y2=0.2025
r6 42 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.2790 $Y=0.2025 $X2=1.2815 $Y2=0.2025
r7 4 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.4040 $Y=0.2025
+ $X2=1.4040 $Y2=0.2340
r8 2 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.2960 $Y=0.2025
+ $X2=1.2960 $Y2=0.2340
r9 38 39 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.4040
+ $Y=0.2340 $X2=1.4175 $Y2=0.2340
r10 37 38 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.3500
+ $Y=0.2340 $X2=1.4040 $Y2=0.2340
r11 36 37 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.2960
+ $Y=0.2340 $X2=1.3500 $Y2=0.2340
r12 18 36 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.2845
+ $Y=0.2340 $X2=1.2960 $Y2=0.2340
r13 21 33 0.624487 $w=2.20462e-08 $l=9.8e-09 $layer=M1 $thickness=3.6e-08
+ $X=1.4310 $Y=0.2340 $X2=1.4310 $Y2=0.2242
r14 21 39 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.4310 $Y=0.2340 $X2=1.4175 $Y2=0.2340
r15 14 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.3895 $Y=0.0675 $X2=1.4020 $Y2=0.0675
r16 35 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.3870 $Y=0.0675 $X2=1.3895 $Y2=0.0675
r17 32 33 0.291487 $w=1.3e-08 $l=1.2e-09 $layer=M1 $thickness=3.6e-08 $X=1.4310
+ $Y=0.2230 $X2=1.4310 $Y2=0.2242
r18 32 31 2.73998 $w=1.3e-08 $l=1.18e-08 $layer=M1 $thickness=3.6e-08 $X=1.4310
+ $Y=0.2230 $X2=1.4310 $Y2=0.2112
r19 30 31 15.4488 $w=1.3e-08 $l=6.62e-08 $layer=M1 $thickness=3.6e-08 $X=1.4310
+ $Y=0.1450 $X2=1.4310 $Y2=0.2112
r20 19 20 5.69636 $w=1.58e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.4310 $Y=0.0675 $X2=1.4310 $Y2=0.0360
r21 19 30 18.0722 $w=1.3e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=1.4310
+ $Y=0.0675 $X2=1.4310 $Y2=0.1450
r22 3 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.4040 $Y=0.0675
+ $X2=1.4040 $Y2=0.0360
r23 20 29 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.4310 $Y=0.0360 $X2=1.4175 $Y2=0.0360
r24 28 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.4040
+ $Y=0.0360 $X2=1.4175 $Y2=0.0360
r25 27 28 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.3500
+ $Y=0.0360 $X2=1.4040 $Y2=0.0360
r26 26 27 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.2960
+ $Y=0.0360 $X2=1.3500 $Y2=0.0360
r27 17 26 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.2845
+ $Y=0.0360 $X2=1.2960 $Y2=0.0360
r28 1 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.2960 $Y=0.0675
+ $X2=1.2960 $Y2=0.0360
r29 25 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.3130 $Y=0.0675 $X2=1.3105 $Y2=0.0675
r30 1 23 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.2960 $Y=0.0675 $X2=1.3105 $Y2=0.0675
r31 13 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.2815 $Y=0.0675 $X2=1.2960 $Y2=0.0675
r32 24 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.2790 $Y=0.0675 $X2=1.2815 $Y2=0.0675
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%CLK VSS 13 3 4 6 1 5
c1 1 VSS 0.00303076f
c2 3 VSS 0.0599481f
c3 4 VSS 0.00256414f
c4 5 VSS 0.00483303f
c5 6 VSS 0.00193917f
r1 5 16 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0630 $X2=0.1080 $Y2=0.0900
r2 15 16 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.0900 $X2=0.1080 $Y2=0.0900
r3 6 9 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0900 $X2=0.0810 $Y2=0.1100
r4 6 15 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0900 $X2=0.0945 $Y2=0.0900
r5 13 12 2.73998 $w=1.3e-08 $l=1.18e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1900 $X2=0.0810 $Y2=0.1782
r6 11 12 3.20636 $w=1.3e-08 $l=1.37e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1645 $X2=0.0810 $Y2=0.1782
r7 10 11 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1530 $X2=0.0810 $Y2=0.1645
r8 8 10 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1530
r9 4 8 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1235 $X2=0.0810 $Y2=0.1350
r10 4 9 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1235 $X2=0.0810 $Y2=0.1100
r11 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r12 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%PD3 VSS 2 4 1
c1 1 VSS 0.000911192f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.0405 $X2=0.7065 $Y2=0.0405
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.0405 $X2=0.6895 $Y2=0.0405
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6895 $Y=0.0405 $X2=0.7065 $Y2=0.0405
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%PD4 VSS 2 4 1
c1 1 VSS 0.00102981f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9890 $Y=0.2295 $X2=0.9765 $Y2=0.2295
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9550 $Y=0.2295 $X2=0.9595 $Y2=0.2295
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9595 $Y=0.2295 $X2=0.9765 $Y2=0.2295
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%noxref_26 VSS 1
c1 1 VSS 0.00433734f
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%PD2 VSS 7 12 4 5 1
c1 1 VSS 0.0074264f
c2 4 VSS 0.00184293f
c3 5 VSS 0.00234071f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7040 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r3 9 5 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.6765
+ $Y=0.2295 $X2=0.7020 $Y2=0.2295
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.6615
+ $Y=0.2295 $X2=0.6765 $Y2=0.2295
r5 1 8 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.6480
+ $Y=0.2295 $X2=0.6615 $Y2=0.2295
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.2295 $X2=0.6460 $Y2=0.2295
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.2295 $X2=0.6335 $Y2=0.2295
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%noxref_27 VSS 1
c1 1 VSS 0.00429939f
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%PD5 VSS 7 12 4 1 5
c1 1 VSS 0.0074251f
c2 4 VSS 0.00187937f
c3 5 VSS 0.00237034f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9890 $Y=0.0405 $X2=0.9865 $Y2=0.0405
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9740 $Y=0.0405 $X2=0.9865 $Y2=0.0405
r3 9 5 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.9585
+ $Y=0.0405 $X2=0.9720 $Y2=0.0405
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.9435
+ $Y=0.0405 $X2=0.9585 $Y2=0.0405
r5 1 8 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.9180
+ $Y=0.0405 $X2=0.9435 $Y2=0.0405
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9035 $Y=0.0405 $X2=0.9160 $Y2=0.0405
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9010 $Y=0.0405 $X2=0.9035 $Y2=0.0405
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%noxref_28 VSS 1
c1 1 VSS 0.00581836f
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%noxref_29 VSS 1
c1 1 VSS 0.00590528f
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%noxref_30 VSS 1
c1 1 VSS 0.0127135f
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%NET13 VSS 12 13 29 8 9 2 7 1
c1 1 VSS 0.00351694f
c2 2 VSS 0.0038088f
c3 7 VSS 0.00294145f
c4 8 VSS 0.0022738f
c5 9 VSS 0.00243954f
r1 29 28 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.0675 $X2=0.6085 $Y2=0.0675
r2 27 28 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6040 $Y=0.0675 $X2=0.6085 $Y2=0.0675
r3 8 27 0.123457 $w=8.1e-08 $l=1e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.0675 $X2=0.6040 $Y2=0.0675
r4 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0675
+ $X2=0.5900 $Y2=0.0720
r5 23 24 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.5805
+ $Y=0.0720 $X2=0.5900 $Y2=0.0720
r6 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0720 $X2=0.5805 $Y2=0.0720
r7 21 22 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.0720 $X2=0.5670 $Y2=0.0720
r8 20 21 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0720 $X2=0.5400 $Y2=0.0720
r9 19 20 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5020
+ $Y=0.0720 $X2=0.5130 $Y2=0.0720
r10 18 19 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4805
+ $Y=0.0720 $X2=0.5020 $Y2=0.0720
r11 17 18 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.4540
+ $Y=0.0720 $X2=0.4805 $Y2=0.0720
r12 16 17 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4440
+ $Y=0.0720 $X2=0.4540 $Y2=0.0720
r13 15 16 1.63233 $w=1.3e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.4370
+ $Y=0.0720 $X2=0.4440 $Y2=0.0720
r14 14 15 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4280
+ $Y=0.0720 $X2=0.4370 $Y2=0.0720
r15 9 14 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4205
+ $Y=0.0720 $X2=0.4280 $Y2=0.0720
r16 1 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4280 $Y2=0.0720
r17 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r18 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r19 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0675 $X2=0.4320 $Y2=0.0675
r20 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4175 $Y2=0.0675
r21 2 8 1e-05
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%MS VSS 10 43 46 50 52 13 17 19 18 3 15 12 1 11 4
+ 14 16
c1 1 VSS 0.00317548f
c2 3 VSS 0.00574996f
c3 4 VSS 0.00955846f
c4 10 VSS 0.0376964f
c5 11 VSS 0.00329686f
c6 12 VSS 0.0031284f
c7 13 VSS 0.00263859f
c8 14 VSS 0.000855829f
c9 15 VSS 0.00355255f
c10 16 VSS 0.00188618f
c11 17 VSS 0.0011264f
c12 18 VSS 0.00137254f
c13 19 VSS 0.00117271f
c14 20 VSS 0.00294923f
r1 52 51 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8810 $Y=0.2295 $X2=0.8785 $Y2=0.2295
r2 13 51 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8660 $Y=0.2295 $X2=0.8785 $Y2=0.2295
r3 12 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.2295 $X2=0.8080 $Y2=0.2295
r4 50 12 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.2295 $X2=0.7955 $Y2=0.2295
r5 47 13 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8370 $Y=0.2295 $X2=0.8640 $Y2=0.2295
r6 4 47 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08 $X=0.8100
+ $Y=0.2295 $X2=0.8370 $Y2=0.2295
r7 4 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8100 $Y=0.2295
+ $X2=0.8100 $Y2=0.2340
r8 15 20 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.2340 $X2=0.8370 $Y2=0.2340
r9 46 45 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8270 $Y=0.0405 $X2=0.8245 $Y2=0.0405
r10 44 45 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8200 $Y=0.0405 $X2=0.8245 $Y2=0.0405
r11 3 44 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8080 $Y=0.0405 $X2=0.8200 $Y2=0.0405
r12 11 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.0405 $X2=0.8080 $Y2=0.0405
r13 43 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.0405 $X2=0.7955 $Y2=0.0405
r14 20 39 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.2340 $X2=0.8370 $Y2=0.2160
r15 3 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8100 $Y=0.0405
+ $X2=0.8100 $Y2=0.0535
r16 38 39 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1870 $X2=0.8370 $Y2=0.2160
r17 37 38 4.89699 $w=1.3e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1660 $X2=0.8370 $Y2=0.1870
r18 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1525 $X2=0.8370 $Y2=0.1660
r19 35 36 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1310 $X2=0.8370 $Y2=0.1525
r20 34 35 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1115 $X2=0.8370 $Y2=0.1310
r21 17 31 1.15159 $w=1.75e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1000 $X2=0.8370 $Y2=0.0900
r22 17 34 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1000 $X2=0.8370 $Y2=0.1115
r23 16 32 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0625 $X2=0.8100 $Y2=0.0720
r24 16 33 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0625 $X2=0.8100 $Y2=0.0535
r25 30 31 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8235 $Y=0.0900 $X2=0.8370 $Y2=0.0900
r26 19 28 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.0900 $X2=0.7965 $Y2=0.0900
r27 19 30 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.0900 $X2=0.8235 $Y2=0.0900
r28 19 32 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0900 $X2=0.8100 $Y2=0.0720
r29 27 28 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.7740
+ $Y=0.0900 $X2=0.7965 $Y2=0.0900
r30 14 27 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7470
+ $Y=0.0900 $X2=0.7740 $Y2=0.0900
r31 14 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7470 $Y=0.0900
+ $X2=0.7500 $Y2=0.0900
r32 14 18 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7470
+ $Y=0.0900 $X2=0.7290 $Y2=0.0900
r33 25 26 5.02115 $w=1.53e-08 $l=8.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.7415 $Y=0.0900 $X2=0.7500 $Y2=0.0900
r34 23 25 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.7385 $Y=0.0900 $X2=0.7415 $Y2=0.0900
r35 1 23 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.7285
+ $Y=0.0900 $X2=0.7385 $Y2=0.0900
r36 1 22 2.48102 $w=2.2e-08 $l=5e-10 $layer=LIG $thickness=4.8e-08 $X=0.7285
+ $Y=0.0900 $X2=0.7290 $Y2=0.0900
r37 22 25 1.47681 $w=1.53e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7290 $Y=0.0900 $X2=0.7415 $Y2=0.0900
r38 10 22 0.314665 $w=2.27e-07 $l=4.5e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.7290 $Y=0.1350 $X2=0.7290 $Y2=0.0900
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%SS VSS 9 34 39 14 13 12 17 16 3 4 15 1 10 11
c1 1 VSS 0.00111166f
c2 3 VSS 0.00569183f
c3 4 VSS 0.00656427f
c4 9 VSS 0.0384074f
c5 10 VSS 0.00326477f
c6 11 VSS 0.00331346f
c7 12 VSS 0.000996827f
c8 13 VSS 0.0084594f
c9 14 VSS 0.00182991f
c10 15 VSS 0.00251753f
c11 16 VSS 0.00670716f
c12 17 VSS 0.00230509f
r1 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0655 $Y=0.2295 $X2=1.0780 $Y2=0.2295
r2 39 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0630 $Y=0.2295 $X2=1.0655 $Y2=0.2295
r3 4 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0800 $Y=0.2295
+ $X2=1.0800 $Y2=0.2340
r4 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.0800
+ $Y=0.2340 $X2=1.0935 $Y2=0.2340
r5 16 32 7.21452 $w=1.425e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.2340 $X2=1.1070 $Y2=0.1980
r6 16 37 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1070 $Y=0.2340 $X2=1.0935 $Y2=0.2340
r7 10 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.0655 $Y=0.0405 $X2=1.0780 $Y2=0.0405
r8 34 10 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.0630 $Y=0.0405 $X2=1.0655 $Y2=0.0405
r9 31 32 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.1440 $X2=1.1070 $Y2=0.1980
r10 14 30 8.95608 $w=1.36627e-08 $l=4.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1070 $Y=0.0810 $X2=1.1070 $Y2=0.0395
r11 14 31 14.691 $w=1.3e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.0810 $X2=1.1070 $Y2=0.1440
r12 3 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0800 $Y=0.0405
+ $X2=1.0800 $Y2=0.0360
r13 17 29 1.40651 $w=1.51875e-08 $l=1.45774e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1070 $Y=0.0305 $X2=1.0935 $Y2=0.0360
r14 17 30 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.0305 $X2=1.1070 $Y2=0.0395
r15 28 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.0800
+ $Y=0.0360 $X2=1.0935 $Y2=0.0360
r16 27 28 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.0685
+ $Y=0.0360 $X2=1.0800 $Y2=0.0360
r17 26 27 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.0640
+ $Y=0.0360 $X2=1.0685 $Y2=0.0360
r18 25 26 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.0360 $X2=1.0640 $Y2=0.0360
r19 13 15 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0260 $Y=0.0360 $X2=0.9990 $Y2=0.0360
r20 13 25 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.0360 $X2=1.0530 $Y2=0.0360
r21 12 22 8.04505 $w=1.3e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.9990
+ $Y=0.0705 $X2=0.9990 $Y2=0.1050
r22 12 15 6.39593 $w=1.55565e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9990 $Y=0.0705 $X2=0.9990 $Y2=0.0360
r23 1 19 2.36633 $w=2.3e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.9990
+ $Y=0.1055 $X2=0.9990 $Y2=0.1055
r24 1 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.9990 $Y=0.1055
+ $X2=0.9990 $Y2=0.1050
r25 9 19 0.314665 $w=2.27e-07 $l=2.95e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.9990 $Y=0.1350 $X2=0.9990 $Y2=0.1055
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%MH VSS 9 55 59 62 66 10 20 14 12 16 3 4 18 17 21
+ 1 19 15
c1 1 VSS 0.000217845f
c2 3 VSS 0.00474068f
c3 4 VSS 0.00496458f
c4 9 VSS 0.036165f
c5 10 VSS 0.0022806f
c6 11 VSS 0.000103794f
c7 12 VSS 0.00212101f
c8 13 VSS 7.09591e-20
c9 14 VSS 0.00911264f
c10 15 VSS 0.00776718f
c11 16 VSS 0.00174852f
c12 17 VSS 0.000662499f
c13 18 VSS 0.000951534f
c14 19 VSS 0.00298815f
c15 20 VSS 5.95945e-20
c16 21 VSS 0.002693f
r1 66 65 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.2295 $X2=0.6085 $Y2=0.2295
r2 64 65 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6040 $Y=0.2295 $X2=0.6085 $Y2=0.2295
r3 3 64 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5920 $Y=0.2295 $X2=0.6040 $Y2=0.2295
r4 13 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2295 $X2=0.5920 $Y2=0.2295
r5 60 61 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.1890 $X2=0.5840 $Y2=0.1890
r6 62 60 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.1890 $X2=0.5795 $Y2=0.1890
r7 12 61 0.185185 $w=5.4e-08 $l=1e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.1890 $X2=0.5840 $Y2=0.1890
r8 12 3 0.518519 $w=3.9e-08 $l=4.05494e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.1890 $X2=0.5920 $Y2=0.2295
r9 59 58 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r10 57 58 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6580 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r11 4 57 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6460 $Y=0.0405 $X2=0.6580 $Y2=0.0405
r12 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0405 $X2=0.6460 $Y2=0.0405
r13 10 4 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0810 $X2=0.6460 $Y2=0.0810
r14 55 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.0810 $X2=0.6335 $Y2=0.0810
r15 3 47 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2295
+ $X2=0.5900 $Y2=0.2340
r16 4 41 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.0405
+ $X2=0.6440 $Y2=0.0360
r17 44 45 1.63233 $w=1.3e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.5990
+ $Y=0.2340 $X2=0.6060 $Y2=0.2340
r18 44 47 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5990
+ $Y=0.2340 $X2=0.5900 $Y2=0.2340
r19 43 45 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.6105
+ $Y=0.2340 $X2=0.6060 $Y2=0.2340
r20 42 43 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6305
+ $Y=0.2340 $X2=0.6105 $Y2=0.2340
r21 14 21 4.53042 $w=1.46981e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6665 $Y=0.2340 $X2=0.6930 $Y2=0.2340
r22 14 42 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.6665
+ $Y=0.2340 $X2=0.6305 $Y2=0.2340
r23 15 39 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.6530
+ $Y=0.0360 $X2=0.6705 $Y2=0.0360
r24 15 41 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6530
+ $Y=0.0360 $X2=0.6440 $Y2=0.0360
r25 21 38 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.2340 $X2=0.6930 $Y2=0.2160
r26 19 33 2.43171 $w=1.804e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6930 $Y=0.0360 $X2=0.6930 $Y2=0.0535
r27 19 39 3.59766 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.0360 $X2=0.6705 $Y2=0.0360
r28 37 38 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1980 $X2=0.6930 $Y2=0.2160
r29 36 37 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1800 $X2=0.6930 $Y2=0.1980
r30 35 36 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1680 $X2=0.6930 $Y2=0.1800
r31 34 35 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1590 $X2=0.6930 $Y2=0.1680
r32 17 20 2.43413 $w=1.59032e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6930 $Y=0.1465 $X2=0.6930 $Y2=0.1310
r33 17 34 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1465 $X2=0.6930 $Y2=0.1590
r34 32 33 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.0625 $X2=0.6930 $Y2=0.0535
r35 31 32 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.0720 $X2=0.6930 $Y2=0.0625
r36 30 31 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.0900 $X2=0.6930 $Y2=0.0720
r37 29 30 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1025 $X2=0.6930 $Y2=0.0900
r38 16 20 2.78392 $w=1.56471e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6930 $Y=0.1140 $X2=0.6930 $Y2=0.1310
r39 16 29 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1140 $X2=0.6930 $Y2=0.1025
r40 20 28 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1310 $X2=0.7110 $Y2=0.1310
r41 27 28 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1310 $X2=0.7110 $Y2=0.1310
r42 18 26 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.1310 $X2=0.7830 $Y2=0.1310
r43 18 27 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.1310 $X2=0.7290 $Y2=0.1310
r44 1 23 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.7830
+ $Y=0.1310 $X2=0.7830 $Y2=0.1310
r45 1 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7830 $Y=0.1310
+ $X2=0.7830 $Y2=0.1310
r46 9 23 0.314665 $w=2.27e-07 $l=4e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.7830 $Y=0.1350 $X2=0.7830 $Y2=0.1310
r47 3 12 1e-05
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%SH VSS 11 12 13 14 84 87 89 92 6 15 16 23 17 25
+ 19 18 5 27 22 2 24 1 20 21 26
c1 1 VSS 0.00253658f
c2 2 VSS 0.0152397f
c3 5 VSS 0.0068362f
c4 6 VSS 0.00696847f
c5 11 VSS 0.0387546f
c6 12 VSS 0.0814369f
c7 13 VSS 0.0814124f
c8 14 VSS 0.0810884f
c9 15 VSS 0.00494096f
c10 16 VSS 0.00514882f
c11 17 VSS 0.00889147f
c12 18 VSS 0.00246706f
c13 19 VSS 0.00213215f
c14 20 VSS 0.00208104f
c15 21 VSS 0.00105832f
c16 22 VSS 0.00502042f
c17 23 VSS 0.00725895f
c18 24 VSS 0.00306415f
c19 25 VSS 0.000988535f
c20 26 VSS 0.00121447f
c21 27 VSS 0.00479346f
r1 92 91 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8810 $Y=0.0405 $X2=0.8785 $Y2=0.0405
r2 5 91 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8660 $Y=0.0405 $X2=0.8785 $Y2=0.0405
r3 88 5 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8540 $Y=0.0405 $X2=0.8660 $Y2=0.0405
r4 15 88 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.0405 $X2=0.8540 $Y2=0.0405
r5 89 15 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.0405 $X2=0.8495 $Y2=0.0405
r6 87 86 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9350 $Y=0.2295 $X2=0.9325 $Y2=0.2295
r7 85 86 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9280 $Y=0.2295 $X2=0.9325 $Y2=0.2295
r8 6 85 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9160 $Y=0.2295 $X2=0.9280 $Y2=0.2295
r9 16 6 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9035 $Y=0.2295 $X2=0.9160 $Y2=0.2295
r10 84 16 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9010 $Y=0.2295 $X2=0.9035 $Y2=0.2295
r11 14 75 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=1.3770
+ $Y=0.1350 $X2=1.3770 $Y2=0.1360
r12 13 69 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=1.3230
+ $Y=0.1350 $X2=1.3230 $Y2=0.1360
r13 12 61 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=1.2690 $Y=0.1350 $X2=1.2690 $Y2=0.1360
r14 5 59 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.0405
+ $X2=0.8640 $Y2=0.0360
r15 6 54 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.9180 $Y=0.2295
+ $X2=0.9180 $Y2=0.2340
r16 73 75 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.3645 $Y=0.1360 $X2=1.3770 $Y2=0.1360
r17 72 73 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.3500 $Y=0.1360 $X2=1.3645 $Y2=0.1360
r18 70 72 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.3355 $Y=0.1360 $X2=1.3500 $Y2=0.1360
r19 69 70 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.3230 $Y=0.1360 $X2=1.3355 $Y2=0.1360
r20 67 69 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.3105 $Y=0.1360 $X2=1.3230 $Y2=0.1360
r21 66 67 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.2960 $Y=0.1360 $X2=1.3105 $Y2=0.1360
r22 64 66 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.2815 $Y=0.1360 $X2=1.2960 $Y2=0.1360
r23 62 64 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=1.2785 $Y=0.1360 $X2=1.2815 $Y2=0.1360
r24 61 62 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=1.2690
+ $Y=0.1360 $X2=1.2785 $Y2=0.1360
r25 2 61 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=1.2595
+ $Y=0.1360 $X2=1.2690 $Y2=0.1360
r26 59 60 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.0360 $X2=0.8775 $Y2=0.0360
r27 57 60 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.0360 $X2=0.8775 $Y2=0.0360
r28 56 57 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.9020
+ $Y=0.0360 $X2=0.8910 $Y2=0.0360
r29 17 24 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.9200
+ $Y=0.0360 $X2=0.9450 $Y2=0.0360
r30 17 56 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.9200
+ $Y=0.0360 $X2=0.9020 $Y2=0.0360
r31 54 55 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.2340 $X2=0.9315 $Y2=0.2340
r32 23 55 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.2340 $X2=0.9315 $Y2=0.2340
r33 51 61 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.2690 $Y=0.1445
+ $X2=1.2690 $Y2=0.1360
r34 22 51 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.2690
+ $Y=0.1085 $X2=1.2690 $Y2=0.1445
r35 24 45 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.0360 $X2=0.9450 $Y2=0.0630
r36 19 40 6.50021 $w=1.33448e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.1980 $X2=0.9450 $Y2=0.1690
r37 19 23 7.21452 $w=1.425e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.1980 $X2=0.9450 $Y2=0.2340
r38 49 51 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=1.2690 $Y=0.1530
+ $X2=1.2690 $Y2=0.1445
r39 48 49 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=1.2445
+ $Y=0.1530 $X2=1.2690 $Y2=0.1530
r40 47 48 9.91056 $w=1.3e-08 $l=4.25e-08 $layer=M2 $thickness=3.6e-08 $X=1.2020
+ $Y=0.1530 $X2=1.2445 $Y2=0.1530
r41 46 47 32.0636 $w=1.3e-08 $l=1.375e-07 $layer=M2 $thickness=3.6e-08
+ $X=1.0645 $Y=0.1530 $X2=1.2020 $Y2=0.1530
r42 27 46 27.8662 $w=1.3e-08 $l=1.195e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.9450 $Y=0.1530 $X2=1.0645 $Y2=0.1530
r43 27 41 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.9450 $Y=0.1530 $X2=0.9450
+ $Y2=0.1485
r44 44 45 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.0900 $X2=0.9450 $Y2=0.0630
r45 43 44 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1000 $X2=0.9450 $Y2=0.0900
r46 42 43 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1100 $X2=0.9450 $Y2=0.1000
r47 18 41 3.96423 $w=1.3e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1315 $X2=0.9450 $Y2=0.1485
r48 18 42 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1315 $X2=0.9450 $Y2=0.1100
r49 39 40 0.4592 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1645 $X2=0.9450 $Y2=0.1690
r50 25 39 0.714311 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1575 $X2=0.9450 $Y2=0.1645
r51 25 41 1.50855 $w=1.55e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1575 $X2=0.9450 $Y2=0.1485
r52 25 27 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.9450 $Y=0.1575 $X2=0.9450
+ $Y2=0.1530
r53 38 40 4.4015 $w=1.35e-08 $l=2.78927e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9720 $Y=0.1620 $X2=0.9450 $Y2=0.1690
r54 37 38 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9990
+ $Y=0.1620 $X2=0.9720 $Y2=0.1620
r55 20 26 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0260 $Y=0.1620 $X2=1.0530 $Y2=0.1620
r56 20 37 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.1620 $X2=0.9990 $Y2=0.1620
r57 26 35 0.915974 $w=2.10182e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0530 $Y=0.1620 $X2=1.0530 $Y2=0.1510
r58 34 35 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1400 $X2=1.0530 $Y2=0.1510
r59 21 34 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1250 $X2=1.0530 $Y2=0.1400
r60 1 31 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=1.0530
+ $Y=0.1400 $X2=1.0530 $Y2=0.1400
r61 1 34 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.0530 $Y=0.1400
+ $X2=1.0530 $Y2=0.1400
r62 11 31 0.314665 $w=2.27e-07 $l=5e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.0530 $Y=0.1350 $X2=1.0530 $Y2=0.1400
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%CLKN VSS 13 14 15 72 74 26 7 22 17 16 19 21 1 8
+ 20 18 29 23 24 3 2 28 25 27
c1 1 VSS 0.00148294f
c2 2 VSS 0.000106006f
c3 3 VSS 0.000190149f
c4 7 VSS 0.00768299f
c5 8 VSS 0.00789839f
c6 13 VSS 0.0592766f
c7 14 VSS 0.00448357f
c8 15 VSS 0.00460295f
c9 16 VSS 0.00618128f
c10 17 VSS 0.00606683f
c11 18 VSS 0.00546167f
c12 19 VSS 0.00364421f
c13 20 VSS 0.00510059f
c14 21 VSS 0.00473615f
c15 22 VSS 0.000611178f
c16 23 VSS 0.000112464f
c17 24 VSS 0.000473001f
c18 25 VSS 0.00356536f
c19 26 VSS 0.00164202f
c20 27 VSS 0.00365958f
c21 28 VSS 0.000153433f
c22 29 VSS 0.0234442f
r1 74 73 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r2 17 73 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r3 72 71 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r4 16 71 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r5 8 69 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0550 $Y2=0.2340
r6 7 66 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0550 $Y2=0.0360
r7 68 69 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.2340 $X2=0.0550 $Y2=0.2340
r8 21 68 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0460 $Y2=0.2340
r9 21 27 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0180 $Y2=0.2340
r10 65 66 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.0360 $X2=0.0550 $Y2=0.0360
r11 20 65 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0460 $Y2=0.0360
r12 20 25 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0180 $Y2=0.0360
r13 27 62 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.2340 $X2=0.0180 $Y2=0.2125
r14 25 61 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.0360 $X2=0.0180 $Y2=0.0630
r15 1 56 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1440
r16 13 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r17 19 26 5.19594 $w=1.44151e-08 $l=2.80401e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1810 $X2=0.0165 $Y2=0.1530
r18 19 62 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1810 $X2=0.0180 $Y2=0.2125
r19 60 61 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0900 $X2=0.0180 $Y2=0.0630
r20 18 26 6.0121 $w=1.425e-08 $l=3.15357e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1215 $X2=0.0165 $Y2=0.1530
r21 18 60 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1215 $X2=0.0180 $Y2=0.0900
r22 2 50 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6210 $Y=0.1350
+ $X2=0.6210 $Y2=0.1395
r23 14 2 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1350
r24 22 56 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1235 $X2=0.1350 $Y2=0.1440
r25 53 54 1.90199 $w=1.38333e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.0255 $Y=0.1530 $X2=0.0345 $Y2=0.1530
r26 26 53 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0165
+ $Y=0.1530 $X2=0.0255 $Y2=0.1530
r27 28 50 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1620 $X2=0.6210 $Y2=0.1395
r28 28 41 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.6210 $Y=0.1620 $X2=0.6210
+ $Y2=0.1530
r29 23 50 5.47996 $w=1.3e-08 $l=2.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1160 $X2=0.6210 $Y2=0.1395
r30 48 49 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1530 $X2=0.1595 $Y2=0.1530
r31 48 56 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1350 $Y=0.1530
+ $X2=0.1350 $Y2=0.1440
r32 47 48 11.8927 $w=1.3e-08 $l=5.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.0840
+ $Y=0.1530 $X2=0.1350 $Y2=0.1530
r33 46 47 11.8927 $w=1.3e-08 $l=5.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.0330
+ $Y=0.1530 $X2=0.0840 $Y2=0.1530
r34 46 54 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.0330 $Y=0.1530
+ $X2=0.0345 $Y2=0.1530
r35 44 49 7.81186 $w=1.3e-08 $l=3.35e-08 $layer=M2 $thickness=3.6e-08 $X=0.1930
+ $Y=0.1530 $X2=0.1595 $Y2=0.1530
r36 43 44 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.2740
+ $Y=0.1530 $X2=0.1930 $Y2=0.1530
r37 41 42 15.2739 $w=1.3e-08 $l=6.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1530 $X2=0.6865 $Y2=0.1530
r38 41 50 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.6210 $Y=0.1530 $X2=0.6210
+ $Y2=0.1395
r39 40 41 34.1623 $w=1.3e-08 $l=1.465e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.4745 $Y=0.1530 $X2=0.6210 $Y2=0.1530
r40 40 43 46.7545 $w=1.3e-08 $l=2.005e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.4745 $Y=0.1530 $X2=0.2740 $Y2=0.1530
r41 29 39 18.3054 $w=1.3e-08 $l=7.85e-08 $layer=M2 $thickness=3.6e-08 $X=0.8125
+ $Y=0.1530 $X2=0.8910 $Y2=0.1530
r42 29 42 29.3819 $w=1.3e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.8125
+ $Y=0.1530 $X2=0.6865 $Y2=0.1530
r43 37 39 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.8910 $Y=0.1440
+ $X2=0.8910 $Y2=0.1530
r44 24 37 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1135 $X2=0.8910 $Y2=0.1440
r45 15 3 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.8910
+ $Y=0.1350 $X2=0.8910 $Y2=0.1350
r46 3 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8910 $Y=0.1350
+ $X2=0.8910 $Y2=0.1440
r47 8 17 1e-05
r48 7 16 1e-05
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%D VSS 4 3 1 5
c1 1 VSS 0.00721328f
c2 3 VSS 0.0461977f
c3 4 VSS 0.00467784f
c4 5 VSS 0.00360385f
r1 5 7 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.1080 $X2=0.4050 $Y2=0.1215
r2 4 7 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1215
r3 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r4 4 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%SE VSS 34 5 6 8 7 11 13 9 12 2 1 10
c1 1 VSS 0.00186245f
c2 2 VSS 0.00396618f
c3 5 VSS 0.0426515f
c4 6 VSS 0.0815892f
c5 7 VSS 0.00157754f
c6 8 VSS 0.000273634f
c7 9 VSS 0.00519189f
c8 10 VSS 0.00504655f
c9 11 VSS 0.000212693f
c10 12 VSS 0.0071379f
c11 13 VSS 0.0505416f
r1 1 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
r2 5 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r3 38 39 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2745
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r4 37 38 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2595
+ $Y=0.1350 $X2=0.2745 $Y2=0.1350
r5 36 37 0.699569 $w=1.3e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.1350 $X2=0.2595 $Y2=0.1350
r6 34 8 2.49951 $w=7.46154e-09 $l=1.95256e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.1340 $X2=0.2445 $Y2=0.1350
r7 8 36 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2445
+ $Y=0.1350 $X2=0.2565 $Y2=0.1350
r8 34 11 0.433689 $w=1.8e-08 $l=4.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.1340 $X2=0.2250 $Y2=0.1297
r9 11 32 3.53073 $w=1.4087e-08 $l=1.72e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.1297 $X2=0.2250 $Y2=0.1125
r10 10 28 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.2250 $Y=0.0360 $X2=0.2250
+ $Y2=0.0450
r11 31 32 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0900 $X2=0.2250 $Y2=0.1125
r12 30 31 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0675 $X2=0.2250 $Y2=0.0900
r13 7 30 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0495 $X2=0.2250 $Y2=0.0675
r14 7 28 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.2250 $Y=0.0495 $X2=0.2250
+ $Y2=0.0450
r15 7 10 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.0495 $X2=0.2250 $Y2=0.0360
r16 28 29 14.108 $w=1.3e-08 $l=6.05e-08 $layer=M2 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0450 $X2=0.2855 $Y2=0.0450
r17 26 29 109.716 $w=1.3e-08 $l=4.705e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.7560 $Y=0.0450 $X2=0.2855 $Y2=0.0450
r18 13 24 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=1.1905
+ $Y=0.0450 $X2=1.2150 $Y2=0.0450
r19 13 26 101.321 $w=1.3e-08 $l=4.345e-07 $layer=M2 $thickness=3.6e-08
+ $X=1.1905 $Y=0.0450 $X2=0.7560 $Y2=0.0450
r20 12 24 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=1.2150 $Y=0.0360 $X2=1.2150
+ $Y2=0.0450
r21 20 21 6.41272 $w=1.3e-08 $l=2.75e-08 $layer=M1 $thickness=3.6e-08 $X=1.2150
+ $Y=0.1085 $X2=1.2150 $Y2=0.1360
r22 19 20 8.51143 $w=1.3e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=1.2150
+ $Y=0.0720 $X2=1.2150 $Y2=0.1085
r23 9 19 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.2150
+ $Y=0.0495 $X2=1.2150 $Y2=0.0720
r24 9 12 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.2150 $Y=0.0495 $X2=1.2150 $Y2=0.0360
r25 9 24 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=1.2150 $Y=0.0495 $X2=1.2150
+ $Y2=0.0450
r26 6 2 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=1.2150
+ $Y=0.1350 $X2=1.2150 $Y2=0.1360
r27 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.2150 $Y=0.1360
+ $X2=1.2150 $Y2=0.1360
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%NET62 VSS 12 13 27 28 7 9 1 2 8
c1 1 VSS 0.00532268f
c2 2 VSS 0.00532842f
c3 7 VSS 0.00334343f
c4 8 VSS 0.00336612f
c5 9 VSS 0.00269386f
r1 28 26 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r2 2 26 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r4 27 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r5 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4280 $Y2=0.1980
r6 21 22 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4185
+ $Y=0.1980 $X2=0.4280 $Y2=0.1980
r7 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1980 $X2=0.4185 $Y2=0.1980
r8 19 20 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.3875
+ $Y=0.1980 $X2=0.4050 $Y2=0.1980
r9 18 19 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3695
+ $Y=0.1980 $X2=0.3875 $Y2=0.1980
r10 17 18 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1980 $X2=0.3695 $Y2=0.1980
r11 16 17 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.1980 $X2=0.3510 $Y2=0.1980
r12 15 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1980 $X2=0.3375 $Y2=0.1980
r13 14 15 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3130
+ $Y=0.1980 $X2=0.3240 $Y2=0.1980
r14 9 14 0.699569 $w=1.3e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.3100
+ $Y=0.1980 $X2=0.3130 $Y2=0.1980
r15 1 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.1980
r16 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r17 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r18 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r19 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%SI VSS 14 3 5 1 4 7 6
c1 1 VSS 0.00582996f
c2 3 VSS 0.00733764f
c3 4 VSS 0.00312402f
c4 5 VSS 0.00302516f
c5 6 VSS 0.00358117f
c6 7 VSS 0.00368725f
r1 6 19 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1980 $X2=0.5130 $Y2=0.1765
r2 5 7 3.2503 $w=1.53684e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1540 $X2=0.5130 $Y2=0.1350
r3 5 19 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1540 $X2=0.5130 $Y2=0.1765
r4 7 16 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1350 $X2=0.4945 $Y2=0.1350
r5 15 16 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4845
+ $Y=0.1350 $X2=0.4945 $Y2=0.1350
r6 14 15 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4750
+ $Y=0.1350 $X2=0.4845 $Y2=0.1350
r7 14 4 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4750
+ $Y=0.1350 $X2=0.4635 $Y2=0.1350
r8 14 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4750 $Y=0.1350
+ $X2=0.4790 $Y2=0.1350
r9 11 12 4.43042 $w=1.53e-08 $l=7.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.4715
+ $Y=0.1350 $X2=0.4790 $Y2=0.1350
r10 9 11 1.86855 $w=1.78125e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.4675 $Y=0.1350 $X2=0.4715 $Y2=0.1350
r11 1 9 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.4575
+ $Y=0.1350 $X2=0.4675 $Y2=0.1350
r12 3 1 2.53453 $w=1.32811e-07 $l=1.5e-09 $layer=LIG $thickness=5.23243e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4575 $Y2=0.1350
r13 3 11 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4715 $Y2=0.1350
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%NET15 VSS 13 24 26 8 1 2 9 11 10
c1 1 VSS 0.00560185f
c2 2 VSS 0.00860417f
c3 8 VSS 0.00326408f
c4 9 VSS 0.00233699f
c5 10 VSS 0.00212701f
c6 11 VSS 0.0210754f
r1 26 25 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r2 10 25 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5420 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r3 9 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4840 $Y2=0.2025
r4 24 9 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r5 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5130 $Y=0.2025
+ $X2=0.4900 $Y2=0.2340
r6 20 21 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4810
+ $Y=0.2340 $X2=0.4900 $Y2=0.2340
r7 19 20 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4690
+ $Y=0.2340 $X2=0.4810 $Y2=0.2340
r8 18 19 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4540
+ $Y=0.2340 $X2=0.4690 $Y2=0.2340
r9 17 18 17.7224 $w=1.3e-08 $l=7.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.4540 $Y2=0.2340
r10 16 17 19.5879 $w=1.3e-08 $l=8.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2940
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r11 15 16 5.59655 $w=1.3e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.2940 $Y2=0.2340
r12 11 15 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2580
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r13 8 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2160
+ $X2=0.2700 $Y2=0.2340
r14 1 8 23.8708 $w=2.02e-08 $l=4.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.2700 $Y=0.1755 $X2=0.2700 $Y2=0.2160
r15 13 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r16 8 12 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r17 2 10 1e-05
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%SEN VSS 9 45 47 16 12 13 4 10 11 14 3 1 15
c1 1 VSS 0.00392544f
c2 3 VSS 0.00838163f
c3 4 VSS 0.00674448f
c4 9 VSS 0.0815978f
c5 10 VSS 0.00418798f
c6 11 VSS 0.00453866f
c7 12 VSS 0.00183276f
c8 13 VSS 0.00367638f
c9 14 VSS 0.000833803f
c10 15 VSS 0.00591401f
c11 16 VSS 0.0158007f
r1 47 46 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.2050 $Y=0.2295 $X2=1.2025 $Y2=0.2295
r2 11 46 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.1900 $Y=0.2295 $X2=1.2025 $Y2=0.2295
r3 4 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.1880 $Y=0.2295
+ $X2=1.1880 $Y2=0.2340
r4 45 44 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.2050 $Y=0.0405 $X2=1.2025 $Y2=0.0405
r5 10 44 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.1900 $Y=0.0405 $X2=1.2025 $Y2=0.0405
r6 41 42 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.1745
+ $Y=0.2340 $X2=1.1880 $Y2=0.2340
r7 15 37 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1610 $Y=0.2340 $X2=1.1610 $Y2=0.2125
r8 15 41 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1610 $Y=0.2340 $X2=1.1745 $Y2=0.2340
r9 39 10 3.98201 $w=3.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.1730 $Y=0.0455 $X2=1.1880 $Y2=0.0455
r10 38 39 3.18561 $w=3.32e-08 $l=1.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.1610 $Y=0.0455 $X2=1.1730 $Y2=0.0455
r11 3 38 3.31834 $w=3.32e-08 $l=1.25e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.1485 $Y=0.0455 $X2=1.1610 $Y2=0.0455
r12 36 37 15.7403 $w=1.3e-08 $l=6.75e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.1450 $X2=1.1610 $Y2=0.2125
r13 35 36 14.9241 $w=1.3e-08 $l=6.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0810 $X2=1.1610 $Y2=0.1450
r14 34 35 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0650 $X2=1.1610 $Y2=0.0810
r15 33 34 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0515 $X2=1.1610 $Y2=0.0650
r16 33 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.1610 $Y=0.0515
+ $X2=1.1610 $Y2=0.0455
r17 32 33 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0425 $X2=1.1610 $Y2=0.0515
r18 13 32 1.28254 $w=1.3e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0370 $X2=1.1610 $Y2=0.0425
r19 30 35 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=1.1610 $Y=0.0810
+ $X2=1.1610 $Y2=0.0810
r20 29 30 27.2832 $w=1.3e-08 $l=1.17e-07 $layer=M2 $thickness=3.6e-08 $X=1.0440
+ $Y=0.0810 $X2=1.1610 $Y2=0.0810
r21 28 29 29.3819 $w=1.3e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.9180
+ $Y=0.0810 $X2=1.0440 $Y2=0.0810
r22 27 28 67.1587 $w=1.3e-08 $l=2.88e-07 $layer=M2 $thickness=3.6e-08 $X=0.6300
+ $Y=0.0810 $X2=0.9180 $Y2=0.0810
r23 26 27 65.0599 $w=1.3e-08 $l=2.79e-07 $layer=M2 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0810 $X2=0.6300 $Y2=0.0810
r24 16 26 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.3395
+ $Y=0.0810 $X2=0.3510 $Y2=0.0810
r25 14 22 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.0720 $X2=0.3510 $Y2=0.0855
r26 14 26 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.3510 $Y=0.0720 $X2=0.3510
+ $Y2=0.0810
r27 22 23 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0855 $X2=0.3510 $Y2=0.0945
r28 22 26 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.3510 $Y=0.0855 $X2=0.3510
+ $Y2=0.0810
r29 21 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1080 $X2=0.3510 $Y2=0.0945
r30 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1215 $X2=0.3510 $Y2=0.1080
r31 12 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1215
r32 9 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r33 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
r34 4 11 1e-05
.ends

.subckt PM_SDFHx3_ASAP7_75t_R%CLKB VSS 14 15 16 17 85 87 26 19 7 18 24 6 20 23
+ 4 22 21 8 2 1 25
c1 1 VSS 0.000273064f
c2 2 VSS 6.64301e-20
c3 3 VSS 1e-36
c4 4 VSS 0.000293845f
c5 6 VSS 0.00737026f
c6 7 VSS 0.00745876f
c7 8 VSS 0.00383969f
c8 14 VSS 0.00581081f
c9 15 VSS 0.00509403f
c10 16 VSS 0.00438215f
c11 17 VSS 0.00521777f
c12 18 VSS 0.00782082f
c13 19 VSS 0.00776725f
c14 20 VSS 0.00337063f
c15 21 VSS 0.00181162f
c16 22 VSS 0.00142377f
c17 23 VSS 0.00610196f
c18 24 VSS 0.00604394f
c19 25 VSS 0.000620286f
c20 26 VSS 0.0245048f
r1 19 7 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1600 $Y2=0.2160
r2 87 19 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r3 18 6 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1600 $Y2=0.0540
r4 85 18 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r5 7 80 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r6 6 77 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r7 1 72 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1355
+ $X2=0.5670 $Y2=0.1350
r8 14 1 3.19489 $w=1.24e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1355
r9 80 81 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r10 24 68 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.1890 $Y2=0.2160
r11 24 81 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2340 $X2=0.1755 $Y2=0.2340
r12 77 78 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r13 23 64 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1890 $Y2=0.0630
r14 23 78 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1755 $Y2=0.0360
r15 25 69 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.1980 $X2=0.5670 $Y2=0.1845
r16 25 54 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.5670 $Y=0.1980 $X2=0.5670
+ $Y2=0.1890
r17 72 73 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1485
r18 70 73 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1620 $X2=0.5670 $Y2=0.1485
r19 21 69 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1755 $X2=0.5670 $Y2=0.1845
r20 21 70 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1755 $X2=0.5670 $Y2=0.1620
r21 67 68 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2035 $X2=0.1890 $Y2=0.2160
r22 66 67 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1990 $X2=0.1890 $Y2=0.2035
r23 65 66 1.28254 $w=1.3e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1935 $X2=0.1890 $Y2=0.1990
r24 63 64 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0900 $X2=0.1890 $Y2=0.0630
r25 62 63 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1100 $X2=0.1890 $Y2=0.0900
r26 61 62 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1325 $X2=0.1890 $Y2=0.1100
r27 60 61 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1540 $X2=0.1890 $Y2=0.1325
r28 59 60 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1655 $X2=0.1890 $Y2=0.1540
r29 58 65 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1845 $X2=0.1890 $Y2=0.1935
r30 20 58 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1735 $X2=0.1890 $Y2=0.1845
r31 20 59 1.86552 $w=1.3e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1735 $X2=0.1890 $Y2=0.1655
r32 55 56 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.6480
+ $Y=0.1890 $X2=0.7290 $Y2=0.1890
r33 54 55 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1890 $X2=0.6480 $Y2=0.1890
r34 54 69 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.5670 $Y=0.1890 $X2=0.5670
+ $Y2=0.1845
r35 53 54 44.0729 $w=1.3e-08 $l=1.89e-07 $layer=M2 $thickness=3.6e-08 $X=0.3780
+ $Y=0.1890 $X2=0.5670 $Y2=0.1890
r36 52 53 44.0729 $w=1.3e-08 $l=1.89e-07 $layer=M2 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1890 $X2=0.3780 $Y2=0.1890
r37 52 58 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1890 $Y=0.1890
+ $X2=0.1890 $Y2=0.1845
r38 26 52 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.1775
+ $Y=0.1890 $X2=0.1890 $Y2=0.1890
r39 4 49 2.78395 $w=2.4e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.9450
+ $Y=0.1780 $X2=0.9450 $Y2=0.1780
r40 17 4 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.9450 $Y=0.1350 $X2=0.9450 $Y2=0.1780
r41 2 42 2.78395 $w=2.4e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.6750
+ $Y=0.1780 $X2=0.6750 $Y2=0.1780
r42 15 2 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.6750 $Y=0.1350 $X2=0.6750 $Y2=0.1780
r43 50 56 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.7290 $Y=0.1845
+ $X2=0.7290 $Y2=0.1890
r44 22 50 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1680 $X2=0.7290 $Y2=0.1845
r45 48 49 6.83711 $w=2.22e-08 $l=1.5e-09 $layer=LISD $thickness=2.7e-08
+ $X=0.9435 $Y=0.1780 $X2=0.9450 $Y2=0.1780
r46 47 48 12.9145 $w=2.22e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9180 $Y=0.1780 $X2=0.9435 $Y2=0.1780
r47 46 47 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9045 $Y=0.1780 $X2=0.9180 $Y2=0.1780
r48 45 46 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8910 $Y=0.1780 $X2=0.9045 $Y2=0.1780
r49 44 45 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8775 $Y=0.1780 $X2=0.8910 $Y2=0.1780
r50 43 44 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8640 $Y=0.1780 $X2=0.8775 $Y2=0.1780
r51 41 42 12.9145 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6885 $Y=0.1780 $X2=0.6750 $Y2=0.1780
r52 40 41 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7155 $Y=0.1780 $X2=0.6885 $Y2=0.1780
r53 38 39 6.07743 $w=2.22e-08 $l=1.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7290 $Y=0.1780 $X2=0.7410 $Y2=0.1780
r54 38 50 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7290 $Y=0.1780
+ $X2=0.7290 $Y2=0.1845
r55 37 38 5.31775 $w=2.22e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7185 $Y=0.1780 $X2=0.7290 $Y2=0.1780
r56 37 40 1.51936 $w=2.22e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.7185
+ $Y=0.1780 $X2=0.7155 $Y2=0.1780
r57 36 39 4.55807 $w=2.22e-08 $l=9e-09 $layer=LISD $thickness=2.7e-08 $X=0.7500
+ $Y=0.1780 $X2=0.7410 $Y2=0.1780
r58 35 36 6.07743 $w=2.22e-08 $l=1.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7620 $Y=0.1780 $X2=0.7500 $Y2=0.1780
r59 34 35 4.05162 $w=2.22e-08 $l=8e-09 $layer=LISD $thickness=2.7e-08 $X=0.7700
+ $Y=0.1780 $X2=0.7620 $Y2=0.1780
r60 33 34 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7835 $Y=0.1780 $X2=0.7700 $Y2=0.1780
r61 32 33 6.58388 $w=2.22e-08 $l=1.3e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7965 $Y=0.1780 $X2=0.7835 $Y2=0.1780
r62 31 32 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8100 $Y=0.1780 $X2=0.7965 $Y2=0.1780
r63 8 31 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8370 $Y=0.1780 $X2=0.8100 $Y2=0.1780
r64 8 43 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8370 $Y=0.1780 $X2=0.8640 $Y2=0.1780
r65 3 30 2.78395 $w=2.4e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.8370
+ $Y=0.1780 $X2=0.8370 $Y2=0.1780
r66 3 8 10.3807 $w=2.30357e-08 $l=0 $layer=LISD $thickness=3.675e-08 $X=0.8370
+ $Y=0.1780 $X2=0.8370 $Y2=0.1780
r67 16 30 0.314665 $w=2.27e-07 $l=4.3e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.8370 $Y=0.1350 $X2=0.8370 $Y2=0.1780
.ends


*
.SUBCKT SDFHx3_ASAP7_75t_R VSS VDD CLK SE D SI QN
*
* VSS VSS
* VDD VDD
* CLK CLK
* SE SE
* D D
* SI SI
* QN QN
*
*

MM20 N_MM20_d N_MM20_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM23 N_MM23_d N_MM22_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM0 N_MM0_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM28 N_MM28_d N_MM2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM29 N_MM29_d N_MM26_g N_MM29_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM27_g N_MM5_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM10_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM6 N_MM6_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM12 N_MM12_d N_MM12_g N_MM12_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM17 N_MM17_d N_MM17_g N_MM17_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM16 N_MM16_d N_MM16_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM14 N_MM14_d N_MM14_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM30 N_MM30_d N_MM30_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM24 N_MM24_d N_MM24_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@3 N_MM24@3_d N_MM24@3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@2 N_MM24@2_d N_MM24@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM21 N_MM21_d N_MM20_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM22 N_MM22_d N_MM22_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g N_MM3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM26 N_MM26_d N_MM26_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM27 N_MM27_d N_MM27_g N_MM27_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM13 N_MM13_d N_MM17_g N_MM13_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM18 N_MM18_d N_MM18_g N_MM18_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM19 N_MM19_d N_MM16_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM15 N_MM15_d N_MM14_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM31 N_MM31_d N_MM30_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM25 N_MM25_d N_MM24_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@3 N_MM25@3_d N_MM24@3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@2 N_MM25@2_d N_MM24@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "SDFHx3_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "SDFHx3_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_SDFHx3_ASAP7_75t_R%NET137 VSS N_MM28_d N_MM29_s N_NET137_1
+ PM_SDFHx3_ASAP7_75t_R%NET137
cc_1 N_NET137_1 N_MM2_g 0.0173478f
cc_2 N_NET137_1 N_MM26_g 0.0172429f
x_PM_SDFHx3_ASAP7_75t_R%noxref_33 VSS N_noxref_33_1
+ PM_SDFHx3_ASAP7_75t_R%noxref_33
cc_3 N_noxref_33_1 N_MM30_g 0.00557982f
cc_4 N_noxref_33_1 N_SEN_3 0.00138104f
cc_5 N_noxref_33_1 N_SEN_10 0.0170354f
cc_6 N_noxref_33_1 N_SS_10 0.000441512f
cc_7 N_noxref_33_1 N_noxref_31_1 0.00768428f
cc_8 N_noxref_33_1 N_noxref_32_1 0.000505958f
x_PM_SDFHx3_ASAP7_75t_R%noxref_34 VSS N_noxref_34_1
+ PM_SDFHx3_ASAP7_75t_R%noxref_34
cc_9 N_noxref_34_1 N_MM30_g 0.00568407f
cc_10 N_noxref_34_1 N_SEN_4 0.000298763f
cc_11 N_noxref_34_1 N_SEN_11 0.0166829f
cc_12 N_noxref_34_1 N_SS_11 0.000611919f
cc_13 N_noxref_34_1 N_noxref_31_1 0.000510566f
cc_14 N_noxref_34_1 N_noxref_32_1 0.00786732f
cc_15 N_noxref_34_1 N_noxref_33_1 0.00152391f
x_PM_SDFHx3_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_SDFHx3_ASAP7_75t_R%noxref_24
cc_16 N_noxref_24_1 N_MM20_g 0.00369504f
cc_17 N_noxref_24_1 N_CLKN_25 5.73325e-20
cc_18 N_noxref_24_1 N_CLKN_26 5.78412e-20
cc_19 N_noxref_24_1 N_CLKN_19 6.38967e-20
cc_20 N_noxref_24_1 N_CLKN_18 0.00031387f
cc_21 N_noxref_24_1 N_CLKN_7 0.000504732f
cc_22 N_noxref_24_1 N_CLKN_16 0.0276256f
x_PM_SDFHx3_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_SDFHx3_ASAP7_75t_R%noxref_25
cc_23 N_noxref_25_1 N_MM20_g 0.00368577f
cc_24 N_noxref_25_1 N_CLKN_27 6.01777e-20
cc_25 N_noxref_25_1 N_CLKN_26 8.78806e-20
cc_26 N_noxref_25_1 N_CLKN_18 0.000151619f
cc_27 N_noxref_25_1 N_CLKN_19 0.000202801f
cc_28 N_noxref_25_1 N_CLKN_8 0.000500585f
cc_29 N_noxref_25_1 N_CLKN_17 0.0276134f
cc_30 N_noxref_25_1 N_noxref_24_1 0.00204371f
x_PM_SDFHx3_ASAP7_75t_R%noxref_31 VSS N_noxref_31_1
+ PM_SDFHx3_ASAP7_75t_R%noxref_31
cc_31 N_noxref_31_1 N_SEN_3 0.00115948f
cc_32 N_noxref_31_1 N_SS_10 0.0170021f
cc_33 N_noxref_31_1 N_MM14_g 0.0057463f
x_PM_SDFHx3_ASAP7_75t_R%noxref_32 VSS N_noxref_32_1
+ PM_SDFHx3_ASAP7_75t_R%noxref_32
cc_34 N_noxref_32_1 N_SEN_11 0.000615803f
cc_35 N_noxref_32_1 N_SS_11 0.0170396f
cc_36 N_noxref_32_1 N_MM14_g 0.00582072f
cc_37 N_noxref_32_1 N_noxref_31_1 0.00153605f
x_PM_SDFHx3_ASAP7_75t_R%NET134 VSS N_MM0_d N_MM5_s N_NET134_7 N_NET134_9
+ N_NET134_1 N_NET134_11 N_NET134_12 N_NET134_10 N_NET134_8 N_NET134_2
+ PM_SDFHx3_ASAP7_75t_R%NET134
cc_38 N_NET134_7 N_SE_1 0.00126947f
cc_39 N_NET134_9 N_SE_10 0.000664316f
cc_40 N_NET134_1 N_SE_8 0.000835188f
cc_41 N_NET134_11 N_SE_7 0.00128985f
cc_42 N_NET134_12 N_SE_10 0.00133731f
cc_43 N_NET134_1 N_MM3_g 0.00158714f
cc_44 N_NET134_11 N_SE_8 0.00366224f
cc_45 N_NET134_10 N_SE_13 0.00425156f
cc_46 N_NET134_7 N_MM3_g 0.0341252f
cc_47 N_NET134_10 N_SEN_12 0.000325017f
cc_48 N_NET134_10 N_SEN_16 0.00037728f
cc_49 N_NET134_11 N_SEN_12 0.00111071f
cc_50 N_NET134_10 N_SEN_14 0.00546661f
cc_51 N_NET134_8 N_SI_1 0.00129807f
cc_52 N_NET134_2 N_MM27_g 0.0015318f
cc_53 N_NET134_8 N_MM27_g 0.0348422f
x_PM_SDFHx3_ASAP7_75t_R%noxref_35 VSS N_noxref_35_1
+ PM_SDFHx3_ASAP7_75t_R%noxref_35
cc_54 N_noxref_35_1 N_MM24@2_g 0.00148629f
cc_55 N_noxref_35_1 N_QN_14 0.0377403f
x_PM_SDFHx3_ASAP7_75t_R%noxref_36 VSS N_noxref_36_1
+ PM_SDFHx3_ASAP7_75t_R%noxref_36
cc_56 N_noxref_36_1 N_MM24@2_g 0.00147703f
cc_57 N_noxref_36_1 N_QN_16 0.0378399f
cc_58 N_noxref_36_1 N_noxref_35_1 0.00177565f
x_PM_SDFHx3_ASAP7_75t_R%QN VSS QN N_MM24_d N_MM24@3_d N_MM24@2_d N_MM25_d
+ N_MM25@3_d N_MM25@2_d N_QN_13 N_QN_19 N_QN_3 N_QN_15 N_QN_4 N_QN_18 N_QN_1
+ N_QN_2 N_QN_16 N_QN_14 PM_SDFHx3_ASAP7_75t_R%QN
cc_59 N_QN_13 N_SH_22 0.00116855f
cc_60 N_QN_13 N_SH_2 0.000442377f
cc_61 N_QN_13 N_MM24@2_g 0.000932857f
cc_62 N_QN_13 N_SH_27 0.000607727f
cc_63 N_QN_19 N_SH_2 0.000816201f
cc_64 N_QN_3 N_MM24@2_g 0.000864538f
cc_65 N_QN_15 N_MM24_g 0.0309949f
cc_66 N_QN_4 N_MM24@2_g 0.000915759f
cc_67 N_QN_18 N_SH_22 0.00122931f
cc_68 N_QN_1 N_MM24_g 0.0021893f
cc_69 N_QN_2 N_SH_22 0.00231951f
cc_70 N_QN_2 N_MM24_g 0.00236173f
cc_71 N_QN_16 N_MM24@2_g 0.0151438f
cc_72 N_QN_15 N_SH_2 0.00690855f
cc_73 N_QN_14 N_MM24@2_g 0.0525879f
cc_74 N_QN_13 N_MM24@3_g 0.0373199f
cc_75 N_QN_13 N_MM24_g 0.0681803f
x_PM_SDFHx3_ASAP7_75t_R%CLK VSS CLK N_MM20_g N_CLK_4 N_CLK_6 N_CLK_1 N_CLK_5
+ PM_SDFHx3_ASAP7_75t_R%CLK
x_PM_SDFHx3_ASAP7_75t_R%PD3 VSS N_MM9_s N_MM8_d N_PD3_1
+ PM_SDFHx3_ASAP7_75t_R%PD3
cc_76 N_PD3_1 N_MM9_g 0.00777391f
cc_77 N_PD3_1 N_MM11_g 0.0078334f
x_PM_SDFHx3_ASAP7_75t_R%PD4 VSS N_MM18_s N_MM19_d N_PD4_1
+ PM_SDFHx3_ASAP7_75t_R%PD4
cc_78 N_PD4_1 N_MM18_g 0.00783221f
cc_79 N_PD4_1 N_MM16_g 0.00773636f
x_PM_SDFHx3_ASAP7_75t_R%noxref_26 VSS N_noxref_26_1
+ PM_SDFHx3_ASAP7_75t_R%noxref_26
cc_80 N_noxref_26_1 N_MM22_g 0.00351361f
cc_81 N_noxref_26_1 N_CLKB_20 0.000144085f
cc_82 N_noxref_26_1 N_CLKB_6 0.00043246f
cc_83 N_noxref_26_1 N_CLKB_18 0.0270419f
cc_84 N_noxref_26_1 N_NET134_7 0.000551932f
x_PM_SDFHx3_ASAP7_75t_R%PD2 VSS N_MM10_s N_MM11_d N_PD2_4 N_PD2_5 N_PD2_1
+ PM_SDFHx3_ASAP7_75t_R%PD2
cc_85 N_PD2_4 N_MM10_g 0.015009f
cc_86 N_PD2_4 N_CLKB_8 0.000126157f
cc_87 N_PD2_4 N_CLKB_2 0.000277575f
cc_88 N_PD2_5 N_CLKB_8 0.0016725f
cc_89 N_PD2_1 N_MM9_g 0.00209556f
cc_90 N_PD2_5 N_MM9_g 0.00734671f
cc_91 N_PD2_4 N_MM9_g 0.0238238f
cc_92 N_PD2_5 N_MM11_g 0.0148543f
cc_93 N_PD2_4 N_MH_14 0.000321607f
cc_94 N_PD2_4 N_MH_3 0.000612749f
cc_95 N_PD2_1 N_MH_14 0.00348597f
x_PM_SDFHx3_ASAP7_75t_R%noxref_27 VSS N_noxref_27_1
+ PM_SDFHx3_ASAP7_75t_R%noxref_27
cc_96 N_noxref_27_1 N_MM22_g 0.00353333f
cc_97 N_noxref_27_1 N_CLKB_20 0.000174169f
cc_98 N_noxref_27_1 N_CLKB_7 0.000434949f
cc_99 N_noxref_27_1 N_CLKB_19 0.026989f
cc_100 N_noxref_27_1 N_NET15_8 0.000588946f
cc_101 N_noxref_27_1 N_noxref_26_1 0.00148613f
x_PM_SDFHx3_ASAP7_75t_R%PD5 VSS N_MM17_s N_MM16_d N_PD5_4 N_PD5_1 N_PD5_5
+ PM_SDFHx3_ASAP7_75t_R%PD5
cc_102 N_PD5_4 N_MM17_g 0.0152561f
cc_103 N_PD5_1 N_MM18_g 0.000757663f
cc_104 N_PD5_5 N_MM18_g 0.00693384f
cc_105 N_PD5_4 N_MM18_g 0.023966f
cc_106 N_PD5_1 N_MM16_g 0.000892138f
cc_107 N_PD5_5 N_MM16_g 0.0156007f
cc_108 N_PD5_1 N_SH_15 0.000514919f
cc_109 N_PD5_1 N_SH_17 0.000490485f
cc_110 N_PD5_1 N_SH_18 0.00057094f
cc_111 N_PD5_4 N_SH_5 0.000658125f
cc_112 N_PD5_1 N_SH_24 0.00237863f
x_PM_SDFHx3_ASAP7_75t_R%noxref_28 VSS N_noxref_28_1
+ PM_SDFHx3_ASAP7_75t_R%noxref_28
cc_113 N_noxref_28_1 N_MM3_g 0.00162919f
cc_114 N_noxref_28_1 N_CLKB_6 9.95779e-20
cc_115 N_noxref_28_1 N_CLKB_18 0.0005185f
cc_116 N_noxref_28_1 N_NET134_7 0.0359613f
cc_117 N_noxref_28_1 N_noxref_26_1 0.00769511f
cc_118 N_noxref_28_1 N_noxref_27_1 0.00046973f
x_PM_SDFHx3_ASAP7_75t_R%noxref_29 VSS N_noxref_29_1
+ PM_SDFHx3_ASAP7_75t_R%noxref_29
cc_119 N_noxref_29_1 N_MM3_g 0.00148085f
cc_120 N_noxref_29_1 N_CLKB_20 0.000107429f
cc_121 N_noxref_29_1 N_CLKB_19 0.00057737f
cc_122 N_noxref_29_1 N_NET15_8 0.0359747f
cc_123 N_noxref_29_1 N_noxref_26_1 0.000466527f
cc_124 N_noxref_29_1 N_noxref_27_1 0.00771769f
cc_125 N_noxref_29_1 N_noxref_28_1 0.00123961f
x_PM_SDFHx3_ASAP7_75t_R%noxref_30 VSS N_noxref_30_1
+ PM_SDFHx3_ASAP7_75t_R%noxref_30
cc_126 N_noxref_30_1 N_MM27_g 0.00149574f
cc_127 N_noxref_30_1 N_SI_1 0.00244779f
cc_128 N_noxref_30_1 N_CLKB_1 0.000186172f
cc_129 N_noxref_30_1 N_MM1_g 0.0107986f
cc_130 N_noxref_30_1 N_NET15_2 0.00115633f
cc_131 N_noxref_30_1 N_NET15_10 0.0161461f
cc_132 N_noxref_30_1 N_NET15_9 0.0551697f
cc_133 N_noxref_30_1 N_NET134_8 0.0370693f
x_PM_SDFHx3_ASAP7_75t_R%NET13 VSS N_MM29_d N_MM5_d N_MM4_s N_NET13_8 N_NET13_9
+ N_NET13_2 N_NET13_7 N_NET13_1 PM_SDFHx3_ASAP7_75t_R%NET13
cc_134 N_NET13_8 N_CLKN_2 0.000897531f
cc_135 N_NET13_9 N_CLKN_23 0.000742582f
cc_136 N_NET13_2 N_MM10_g 0.000866178f
cc_137 N_NET13_9 N_CLKN_29 0.00092171f
cc_138 N_NET13_8 N_MM10_g 0.0327369f
cc_139 N_NET13_9 N_SE_13 0.00227277f
cc_140 N_NET13_9 N_MM2_g 0.000309987f
cc_141 N_NET13_9 N_SEN_12 0.000111384f
cc_142 N_NET13_9 N_SEN_14 0.000544157f
cc_143 N_NET13_9 N_SEN_16 0.00391645f
cc_144 N_NET13_7 N_D_1 0.000880873f
cc_145 N_NET13_1 N_MM26_g 0.00126271f
cc_146 N_NET13_9 N_D_5 0.0027194f
cc_147 N_NET13_7 N_MM26_g 0.0342508f
cc_148 N_NET13_9 N_SI_4 0.000432229f
cc_149 N_NET13_1 N_MM27_g 0.000757232f
cc_150 N_NET13_7 N_SI_1 0.00082035f
cc_151 N_NET13_9 N_SI_7 0.00250552f
cc_152 N_NET13_7 N_MM27_g 0.0334618f
cc_153 N_NET13_8 N_CLKB_21 0.000153116f
cc_154 N_NET13_8 N_CLKB_1 0.00110832f
cc_155 N_NET13_2 N_MM1_g 0.00116654f
cc_156 N_NET13_9 N_CLKB_21 0.00236413f
cc_157 N_NET13_8 N_MM1_g 0.0355738f
cc_158 N_NET13_8 N_MH_10 0.00114778f
cc_159 N_NET13_9 N_MH_15 0.000948505f
cc_160 N_NET13_2 N_MH_4 0.00367665f
cc_161 N_NET13_7 N_NET134_10 0.000583242f
cc_162 N_NET13_9 N_NET134_2 0.000634232f
cc_163 N_NET13_7 N_NET134_8 0.000642297f
cc_164 N_NET13_1 N_NET134_2 0.00381259f
cc_165 N_NET13_9 N_NET134_10 0.00907183f
x_PM_SDFHx3_ASAP7_75t_R%MS VSS N_MM11_g N_MM6_d N_MM12_d N_MM7_d N_MM13_d
+ N_MS_13 N_MS_17 N_MS_19 N_MS_18 N_MS_3 N_MS_15 N_MS_12 N_MS_1 N_MS_11 N_MS_4
+ N_MS_14 N_MS_16 PM_SDFHx3_ASAP7_75t_R%MS
cc_166 N_MS_13 N_CLKN_24 0.000245511f
cc_167 N_MS_13 N_MM10_g 0.000137844f
cc_168 N_MS_13 N_CLKN_29 0.000349468f
cc_169 N_MS_13 N_CLKN_3 0.000222252f
cc_170 N_MS_17 N_CLKN_24 0.0045445f
cc_171 N_MS_17 N_CLKN_3 0.000289706f
cc_172 N_MS_19 N_CLKN_24 0.000418989f
cc_173 N_MS_18 N_CLKN_29 0.0016246f
cc_174 N_MS_13 N_MM17_g 0.0155046f
cc_175 N_MS_18 N_SEN_16 0.00092503f
cc_176 N_MS_19 N_SEN_16 0.0030369f
cc_177 N_MS_3 N_CLKB_22 0.00014273f
cc_178 N_MS_3 N_CLKB_8 0.000652432f
cc_179 N_MS_3 N_CLKB_2 9.25654e-20
cc_180 N_MS_3 N_CLKB_26 0.000142007f
cc_181 N_MS_15 N_CLKB_22 0.000281055f
cc_182 N_MS_13 N_MM12_g 0.00786932f
cc_183 N_MS_15 N_CLKB_8 0.000361999f
cc_184 N_MS_12 N_MM12_g 0.00781547f
cc_185 N_MS_1 N_MM9_g 0.000704144f
cc_186 N_MS_17 N_CLKB_8 0.00154178f
cc_187 N_MS_11 N_MM12_g 0.006509f
cc_188 N_MS_4 N_MM12_g 0.00257216f
cc_189 N_MS_4 N_CLKB_8 0.00639207f
cc_190 N_MM11_g N_MM9_g 0.0141709f
cc_191 N_MS_3 N_MM12_g 0.0259821f
x_PM_SDFHx3_ASAP7_75t_R%SS VSS N_MM16_g N_MM14_d N_MM15_d N_SS_14 N_SS_13
+ N_SS_12 N_SS_17 N_SS_16 N_SS_3 N_SS_4 N_SS_15 N_SS_1 N_SS_10 N_SS_11
+ PM_SDFHx3_ASAP7_75t_R%SS
cc_192 N_SS_14 N_SE_13 0.000528394f
cc_193 N_SS_13 N_SE_13 0.000906364f
cc_194 N_SS_12 N_SE_13 0.00296079f
cc_195 N_SS_14 N_SEN_3 0.00122843f
cc_196 N_SS_14 N_SEN_4 0.000105992f
cc_197 N_SS_14 N_SEN_15 0.000108856f
cc_198 N_SS_13 N_SEN_16 0.00035578f
cc_199 N_SS_17 N_SEN_13 0.000424246f
cc_200 N_SS_16 N_SEN_15 0.000788228f
cc_201 N_SS_12 N_SEN_16 0.00262193f
cc_202 N_SS_14 N_SEN_13 0.00845023f
cc_203 N_MM16_g N_CLKB_8 0.000681165f
cc_204 N_MM16_g N_CLKB_4 0.000426619f
cc_205 N_MM16_g N_MM18_g 0.0133584f
x_PM_SDFHx3_ASAP7_75t_R%MH VSS N_MM7_g N_MM4_d N_MM9_d N_MM1_d N_MM10_d N_MH_10
+ N_MH_20 N_MH_14 N_MH_12 N_MH_16 N_MH_3 N_MH_4 N_MH_18 N_MH_17 N_MH_21 N_MH_1
+ N_MH_19 N_MH_15 PM_SDFHx3_ASAP7_75t_R%MH
cc_206 N_MH_10 N_CLKN_23 0.000252056f
cc_207 N_MH_10 N_CLKN_3 0.00010979f
cc_208 N_MH_10 N_MM17_g 0.000137032f
cc_209 N_MH_10 N_CLKN_28 0.00029397f
cc_210 N_MH_20 N_CLKN_28 0.00031886f
cc_211 N_MH_14 N_CLKN_28 0.000451586f
cc_212 N_MH_12 N_MM10_g 0.0163723f
cc_213 N_MH_16 N_CLKN_23 0.000527215f
cc_214 N_MH_3 N_CLKN_2 0.000605158f
cc_215 N_MH_4 N_CLKN_23 0.000808312f
cc_216 N_MH_18 N_CLKN_29 0.000902915f
cc_217 N_MH_4 N_MM10_g 0.00111142f
cc_218 N_MH_3 N_MM10_g 0.00122492f
cc_219 N_MH_10 N_CLKN_2 0.00160875f
cc_220 N_MH_17 N_CLKN_29 0.00166213f
cc_221 N_MH_17 N_CLKN_28 0.00210986f
cc_222 N_MH_10 N_MM10_g 0.0527099f
cc_223 N_MH_10 N_CLKB_21 0.000122674f
cc_224 N_MH_10 N_CLKB_22 0.000341104f
cc_225 N_MH_10 N_MM1_g 0.000428406f
cc_226 N_MH_10 N_CLKB_1 0.000203064f
cc_227 N_MH_3 N_CLKB_21 0.000340472f
cc_228 N_MH_3 N_CLKB_25 0.000359477f
cc_229 N_MH_21 N_CLKB_22 0.000404124f
cc_230 N_MH_17 N_CLKB_22 0.0064603f
cc_231 N_MH_17 N_CLKB_2 0.000497541f
cc_232 N_MH_1 N_CLKB_8 0.00208585f
cc_233 N_MH_4 N_MM9_g 0.000633766f
cc_234 N_MH_12 N_CLKB_1 0.00066955f
cc_235 N_MH_17 N_CLKB_8 0.000774024f
cc_236 N_MH_14 N_CLKB_26 0.00145898f
cc_237 N_MH_18 N_CLKB_22 0.00150019f
cc_238 N_MH_3 N_MM1_g 0.0015637f
cc_239 N_MH_14 N_CLKB_25 0.00372211f
cc_240 N_MM7_g N_CLKB_8 0.00508685f
cc_241 N_MH_12 N_MM1_g 0.0330064f
cc_242 N_MM7_g N_MM12_g 0.01274f
cc_243 N_MH_10 N_MM9_g 0.0361728f
cc_244 N_MH_19 N_MS_18 0.000267301f
cc_245 N_MH_4 N_MS_1 0.00036046f
cc_246 N_MH_18 N_MS_19 0.000373988f
cc_247 N_MH_18 N_MS_1 0.000662927f
cc_248 N_MM7_g N_MS_3 0.000937847f
cc_249 N_MH_18 N_MS_17 0.000995278f
cc_250 N_MH_1 N_MS_14 0.00100343f
cc_251 N_MH_1 N_MS_1 0.00130262f
cc_252 N_MM7_g N_MS_12 0.00632604f
cc_253 N_MM7_g N_MS_1 0.00241313f
cc_254 N_MM7_g N_MS_11 0.00639585f
cc_255 N_MH_18 N_MS_14 0.0045934f
cc_256 N_MH_16 N_MS_18 0.00497526f
cc_257 N_MM7_g N_MM11_g 0.0294071f
x_PM_SDFHx3_ASAP7_75t_R%SH VSS N_MM14_g N_MM24_g N_MM24@3_g N_MM24@2_g N_MM13_s
+ N_MM18_d N_MM12_s N_MM17_d N_SH_6 N_SH_15 N_SH_16 N_SH_23 N_SH_17 N_SH_25
+ N_SH_19 N_SH_18 N_SH_5 N_SH_27 N_SH_22 N_SH_2 N_SH_24 N_SH_1 N_SH_20 N_SH_21
+ N_SH_26 PM_SDFHx3_ASAP7_75t_R%SH
cc_258 N_SH_6 N_MM17_g 0.000158318f
cc_259 N_SH_15 N_MM17_g 0.00676966f
cc_260 N_SH_16 N_MM17_g 0.00683991f
cc_261 N_SH_23 N_CLKN_24 0.000285603f
cc_262 N_SH_17 N_CLKN_24 0.000369687f
cc_263 N_SH_25 N_CLKN_24 0.000402567f
cc_264 N_SH_19 N_CLKN_24 0.00046657f
cc_265 N_SH_18 N_CLKN_3 0.000570191f
cc_266 N_SH_5 N_CLKN_3 0.000576027f
cc_267 N_SH_27 N_CLKN_29 0.000763609f
cc_268 N_SH_18 N_CLKN_24 0.00451947f
cc_269 N_SH_17 N_CLKN_29 0.0011137f
cc_270 N_SH_5 N_MM17_g 0.0183294f
cc_271 N_SH_22 N_SE_12 0.000230203f
cc_272 N_SH_18 N_SE_13 0.000315749f
cc_273 N_SH_2 N_SE_2 0.00175819f
cc_274 N_SH_17 N_SE_13 0.00102295f
cc_275 N_SH_27 N_SE_13 0.00207802f
cc_276 N_SH_24 N_SE_13 0.00271358f
cc_277 N_MM24_g N_MM30_g 0.00337871f
cc_278 N_SH_22 N_SE_9 0.00615509f
cc_279 N_SH_24 N_SEN_16 4.73311e-20
cc_280 N_MM24_g N_SEN_3 5.1306e-20
cc_281 N_SH_1 N_SEN_13 0.00014553f
cc_282 N_SH_20 N_SEN_16 0.000109197f
cc_283 N_SH_27 N_SEN_15 0.000118258f
cc_284 N_SH_22 N_SEN_13 0.000156473f
cc_285 N_SH_27 N_SEN_13 0.00151323f
cc_286 N_SH_22 N_SEN_15 0.000259176f
cc_287 N_SH_21 N_SEN_16 0.000283404f
cc_288 N_SH_17 N_SEN_16 0.000374992f
cc_289 N_SH_27 N_SEN_16 0.00450355f
cc_290 N_SH_18 N_SEN_16 0.00607529f
cc_291 N_SH_16 N_CLKB_8 8.2715e-20
cc_292 N_SH_16 N_CLKB_26 8.49552e-20
cc_293 N_MM14_g N_MM18_g 8.8363e-20
cc_294 N_SH_23 N_CLKB_8 0.000196954f
cc_295 N_SH_25 N_CLKB_8 0.000203975f
cc_296 N_SH_15 N_MM12_g 0.00680288f
cc_297 N_SH_6 N_CLKB_8 0.000276295f
cc_298 N_SH_20 N_CLKB_8 0.000396208f
cc_299 N_SH_18 N_CLKB_8 0.000448364f
cc_300 N_SH_19 N_CLKB_8 0.000605537f
cc_301 N_SH_16 N_CLKB_4 0.000673075f
cc_302 N_SH_6 N_MM18_g 0.00100239f
cc_303 N_SH_5 N_CLKB_8 0.0028297f
cc_304 N_SH_5 N_MM12_g 0.00948039f
cc_305 N_SH_16 N_MM18_g 0.0160001f
cc_306 N_SH_19 N_MS_3 9.84548e-20
cc_307 N_SH_23 N_MS_3 0.000179155f
cc_308 N_SH_16 N_MS_3 0.000436412f
cc_309 N_SH_6 N_MS_3 0.000220896f
cc_310 N_SH_15 N_MS_3 0.000232021f
cc_311 N_SH_15 N_MS_11 0.000234022f
cc_312 N_SH_23 N_MS_4 0.000335705f
cc_313 N_SH_6 N_MS_4 0.000424812f
cc_314 N_SH_17 N_MS_16 0.00043823f
cc_315 N_SH_23 N_MS_17 0.000517956f
cc_316 N_SH_16 N_MS_4 0.00059315f
cc_317 N_SH_17 N_MS_19 0.00132439f
cc_318 N_SH_5 N_MS_3 0.00373295f
cc_319 N_SH_19 N_MM16_g 9.92316e-20
cc_320 N_SH_21 N_SS_13 0.000311072f
cc_321 N_MM14_g N_SS_3 0.000322901f
cc_322 N_MM14_g N_SS_4 0.00042065f
cc_323 N_SH_24 N_SS_15 0.000580125f
cc_324 N_SH_26 N_SS_16 0.000641443f
cc_325 N_SH_26 N_SS_14 0.00069774f
cc_326 N_SH_18 N_SS_1 0.000810777f
cc_327 N_SH_1 N_SS_14 0.000948913f
cc_328 N_MM14_g N_SS_1 0.00111318f
cc_329 N_SH_1 N_MM16_g 0.00135492f
cc_330 N_SH_20 N_SS_12 0.00154855f
cc_331 N_SH_27 N_SS_14 0.00174157f
cc_332 N_MM14_g N_SS_10 0.00649586f
cc_333 N_MM14_g N_SS_11 0.00660051f
cc_334 N_SH_18 N_SS_12 0.00462671f
cc_335 N_SH_21 N_SS_14 0.00485052f
cc_336 N_MM14_g N_MM16_g 0.0300227f
x_PM_SDFHx3_ASAP7_75t_R%CLKN VSS N_MM22_g N_MM10_g N_MM17_g N_MM20_d N_MM21_d
+ N_CLKN_26 N_CLKN_7 N_CLKN_22 N_CLKN_17 N_CLKN_16 N_CLKN_19 N_CLKN_21 N_CLKN_1
+ N_CLKN_8 N_CLKN_20 N_CLKN_18 N_CLKN_29 N_CLKN_23 N_CLKN_24 N_CLKN_3 N_CLKN_2
+ N_CLKN_28 N_CLKN_25 N_CLKN_27 PM_SDFHx3_ASAP7_75t_R%CLKN
cc_337 N_CLKN_26 N_MM20_g 0.000235607f
cc_338 N_CLKN_7 N_MM20_g 0.00109794f
cc_339 N_CLKN_22 N_MM20_g 0.000270134f
cc_340 N_CLKN_17 N_MM20_g 0.011216f
cc_341 N_CLKN_16 N_MM20_g 0.011219f
cc_342 N_CLKN_19 N_CLK_4 0.000469867f
cc_343 N_CLKN_21 N_CLK_4 0.000484622f
cc_344 N_CLKN_1 N_CLK_6 0.000644362f
cc_345 N_CLKN_8 N_MM20_g 0.000752868f
cc_346 N_CLKN_26 N_CLK_1 0.000930979f
cc_347 N_CLKN_20 N_CLK_6 0.000991634f
cc_348 N_CLKN_22 N_CLK_6 0.00104499f
cc_349 N_CLKN_18 N_CLK_6 0.00109768f
cc_350 N_CLKN_29 N_CLK_6 0.00129286f
cc_351 N_CLKN_22 N_CLK_4 0.00147124f
cc_352 N_CLKN_20 N_CLK_5 0.00188064f
cc_353 N_CLKN_1 N_CLK_1 0.002428f
cc_354 N_CLKN_26 N_CLK_4 0.00645141f
cc_355 N_MM22_g N_MM20_g 0.0351946f
x_PM_SDFHx3_ASAP7_75t_R%D VSS D N_MM26_g N_D_1 N_D_5 PM_SDFHx3_ASAP7_75t_R%D
cc_356 N_MM26_g N_SEN_16 0.000472395f
cc_357 N_MM26_g N_SEN_1 0.000865616f
cc_358 N_D_1 N_SEN_1 0.00120732f
cc_359 N_D_5 N_SEN_14 0.0015929f
cc_360 N_D N_SEN_12 0.00215936f
cc_361 N_MM26_g N_MM2_g 0.00504614f
x_PM_SDFHx3_ASAP7_75t_R%SE VSS SE N_MM3_g N_MM30_g N_SE_8 N_SE_7 N_SE_11
+ N_SE_13 N_SE_9 N_SE_12 N_SE_2 N_SE_1 N_SE_10 PM_SDFHx3_ASAP7_75t_R%SE
cc_362 N_SE_8 N_CLKN_23 3.39836e-20
cc_363 N_SE_7 N_CLKN_18 3.51048e-20
cc_364 N_SE_11 N_CLKN_1 3.66514e-20
cc_365 N_SE_11 N_CLKN_22 5.50724e-20
cc_366 N_SE_7 N_CLKN_29 0.000403674f
cc_367 N_SE_11 N_CLKN_29 0.000313663f
cc_368 N_SE_13 N_CLKN_24 0.00050805f
cc_369 N_SE_13 N_CLKN_29 0.00246287f
cc_370 N_SE_8 N_CLKN_29 0.00356891f
x_PM_SDFHx3_ASAP7_75t_R%NET62 VSS N_MM3_s N_MM2_d N_MM26_d N_MM27_s N_NET62_7
+ N_NET62_9 N_NET62_1 N_NET62_2 N_NET62_8 PM_SDFHx3_ASAP7_75t_R%NET62
cc_371 N_NET62_7 N_SE_1 0.00103247f
cc_372 N_NET62_9 N_SE_8 0.000684929f
cc_373 N_NET62_1 N_MM3_g 0.000836295f
cc_374 N_NET62_7 N_MM3_g 0.032969f
cc_375 N_NET62_7 N_SEN_1 0.000921407f
cc_376 N_NET62_1 N_MM2_g 0.000853056f
cc_377 N_NET62_9 N_SEN_12 0.00218916f
cc_378 N_NET62_7 N_MM2_g 0.0330302f
cc_379 N_NET62_2 N_MM26_g 0.000866372f
cc_380 N_NET62_9 N_D 0.00225396f
cc_381 N_NET62_8 N_MM26_g 0.0340503f
cc_382 N_NET62_9 N_SI_4 0.000662149f
cc_383 N_NET62_8 N_SI_1 0.00077815f
cc_384 N_NET62_2 N_MM27_g 0.000817129f
cc_385 N_NET62_8 N_MM27_g 0.0335868f
cc_386 N_NET62_9 N_CLKB_26 0.00296544f
cc_387 N_NET62_2 N_NET15_11 0.000548255f
cc_388 N_NET62_7 N_NET15_8 0.00110602f
cc_389 N_NET62_8 N_NET15_9 0.000555324f
cc_390 N_NET62_1 N_NET15_11 0.000598084f
cc_391 N_NET62_8 N_NET15_2 0.00130113f
cc_392 N_NET62_2 N_NET15_2 0.00161309f
cc_393 N_NET62_1 N_NET15_1 0.00303285f
cc_394 N_NET62_9 N_NET15_11 0.0130952f
x_PM_SDFHx3_ASAP7_75t_R%SI VSS SI N_MM27_g N_SI_5 N_SI_1 N_SI_4 N_SI_7 N_SI_6
+ PM_SDFHx3_ASAP7_75t_R%SI
cc_395 N_SI_5 N_CLKN_29 0.00248818f
cc_396 N_SI_1 N_MM26_g 0.000900113f
cc_397 N_SI_4 N_D_5 0.00100829f
cc_398 N_MM27_g N_MM26_g 0.00404443f
x_PM_SDFHx3_ASAP7_75t_R%NET15 VSS N_MM3_d N_MM27_d N_MM1_s N_NET15_8 N_NET15_1
+ N_NET15_2 N_NET15_9 N_NET15_11 N_NET15_10 PM_SDFHx3_ASAP7_75t_R%NET15
cc_399 N_NET15_8 N_SE_8 0.000706896f
cc_400 N_NET15_8 N_SE_1 0.00106011f
cc_401 N_NET15_1 N_MM3_g 0.00131293f
cc_402 N_NET15_8 N_MM3_g 0.0340628f
cc_403 N_NET15_2 N_SI_5 0.000638001f
cc_404 N_NET15_9 N_SI_1 0.00143375f
cc_405 N_NET15_2 N_SI_6 0.00293121f
cc_406 N_NET15_11 N_SI_6 0.00308262f
cc_407 N_NET15_9 N_MM27_g 0.0349635f
cc_408 N_NET15_10 N_CLKB_20 4.86963e-20
cc_409 N_NET15_10 N_CLKB_24 0.000286139f
cc_410 N_NET15_10 N_CLKB_7 0.000132828f
cc_411 N_NET15_10 N_CLKB_19 0.000143024f
cc_412 N_NET15_10 N_CLKB_1 0.00102103f
cc_413 N_NET15_10 N_CLKB_25 0.000339884f
cc_414 N_NET15_10 N_CLKB_21 0.000351015f
cc_415 N_NET15_1 N_CLKB_20 0.00092126f
cc_416 N_NET15_2 N_MM1_g 0.00158754f
cc_417 N_NET15_11 N_CLKB_26 0.00363633f
cc_418 N_NET15_10 N_MM1_g 0.0338671f
cc_419 N_NET15_2 N_MH_3 0.00118685f
cc_420 N_NET15_2 N_MH_12 0.00289139f
x_PM_SDFHx3_ASAP7_75t_R%SEN VSS N_MM2_g N_MM30_d N_MM31_d N_SEN_16 N_SEN_12
+ N_SEN_13 N_SEN_4 N_SEN_10 N_SEN_11 N_SEN_14 N_SEN_3 N_SEN_1 N_SEN_15
+ PM_SDFHx3_ASAP7_75t_R%SEN
cc_421 N_SEN_16 N_CLKN_24 0.00295699f
cc_422 N_SEN_16 N_CLKN_23 0.000503602f
cc_423 N_SEN_12 N_CLKN_29 0.00327925f
cc_424 N_SEN_16 N_CLKN_29 0.0107478f
cc_425 N_SEN_13 N_SE_9 0.00782246f
cc_426 N_SEN_4 N_SE_9 0.000213952f
cc_427 N_SEN_10 N_MM30_g 0.0232223f
cc_428 N_SEN_11 N_MM30_g 0.0067982f
cc_429 N_SEN_14 N_SE_13 0.000247294f
cc_430 N_SEN_3 N_SE_9 0.000259952f
cc_431 N_SEN_1 N_SE_8 0.000309112f
cc_432 N_SEN_13 N_SE_12 0.000329572f
cc_433 N_SEN_4 N_MM30_g 0.000355273f
cc_434 N_SEN_3 N_SE_2 0.000413508f
cc_435 N_SEN_15 N_SE_9 0.000417746f
cc_436 N_SEN_1 N_SE_1 0.00129184f
cc_437 N_SEN_13 N_SE_2 0.000422208f
cc_438 N_SEN_12 N_SE_13 0.000479966f
cc_439 N_SEN_13 N_SE_13 0.000514992f
cc_440 N_SEN_3 N_MM30_g 0.000947816f
cc_441 N_SEN_12 N_SE_8 0.00172568f
cc_442 N_MM2_g N_MM3_g 0.00330887f
cc_443 N_SEN_16 N_SE_13 0.0652305f
x_PM_SDFHx3_ASAP7_75t_R%CLKB VSS N_MM1_g N_MM9_g N_MM12_g N_MM18_g N_MM23_d
+ N_MM22_d N_CLKB_26 N_CLKB_19 N_CLKB_7 N_CLKB_18 N_CLKB_24 N_CLKB_6 N_CLKB_20
+ N_CLKB_23 N_CLKB_4 N_CLKB_22 N_CLKB_21 N_CLKB_8 N_CLKB_2 N_CLKB_1 N_CLKB_25
+ PM_SDFHx3_ASAP7_75t_R%CLKB
cc_444 N_CLKB_26 N_CLK_5 5.1445e-20
cc_445 N_CLKB_19 N_CLK_5 7.11297e-20
cc_446 N_CLKB_7 N_CLK_5 0.000491718f
cc_447 N_CLKB_18 N_CLK_5 8.91394e-20
cc_448 N_CLKB_24 N_CLK_5 0.000113024f
cc_449 N_CLKB_6 N_CLK_5 0.000386069f
cc_450 N_CLKB_20 N_CLK_6 0.000427282f
cc_451 N_CLKB_23 N_CLK_5 0.00187738f
cc_452 N_CLKB_23 N_CLKN_29 2.90609e-20
cc_453 N_CLKB_24 N_CLKN_29 3.80829e-20
cc_454 N_CLKB_23 N_CLKN_18 4.19252e-20
cc_455 N_CLKB_6 N_MM22_g 0.000651679f
cc_456 N_CLKB_24 N_CLKN_21 9.37071e-20
cc_457 N_CLKB_7 N_MM22_g 0.000788053f
cc_458 N_CLKB_4 N_MM17_g 0.000208159f
cc_459 N_CLKB_23 N_CLKN_22 0.000268624f
cc_460 N_CLKB_22 N_CLKN_29 0.000676953f
cc_461 N_CLKB_21 N_CLKN_29 0.00032759f
cc_462 N_CLKB_20 N_CLKN_22 0.00454098f
cc_463 N_CLKB_24 N_CLKN_22 0.000383004f
cc_464 N_CLKB_18 N_MM22_g 0.0386421f
cc_465 N_CLKB_19 N_MM22_g 0.0111504f
cc_466 N_CLKB_26 N_CLKN_23 0.000478614f
cc_467 N_CLKB_20 N_CLKN_29 0.00052875f
cc_468 N_CLKB_8 N_CLKN_24 0.000531969f
cc_469 N_CLKB_2 N_MM10_g 0.000560153f
cc_470 N_CLKB_20 N_CLKN_1 0.000579205f
cc_471 N_CLKB_8 N_CLKN_3 0.0027913f
cc_472 N_CLKB_19 N_CLKN_1 0.000784303f
cc_473 N_CLKB_1 N_CLKN_2 0.00223836f
cc_474 N_CLKB_25 N_CLKN_28 0.00165668f
cc_475 N_CLKB_21 N_CLKN_23 0.00265808f
cc_476 N_MM9_g N_MM10_g 0.00370557f
cc_477 N_CLKB_8 N_MM17_g 0.00493104f
cc_478 N_MM18_g N_MM17_g 0.00578286f
cc_479 N_MM1_g N_MM10_g 0.00704327f
cc_480 N_MM12_g N_MM17_g 0.0182761f
cc_481 N_CLKB_26 N_CLKN_29 0.0458181f
cc_482 N_CLKB_7 N_SE_11 4.71947e-20
cc_483 N_CLKB_6 N_SE_11 5.44479e-20
cc_484 N_MM18_g N_SE_13 0.000107802f
cc_485 N_CLKB_6 N_SE_7 0.000174715f
cc_486 N_CLKB_26 N_SE_13 0.000265f
cc_487 N_CLKB_23 N_SE_7 0.000351201f
cc_488 N_CLKB_21 N_SE_13 0.000837093f
cc_489 N_CLKB_26 N_SE_8 0.00121501f
cc_490 N_CLKB_23 N_SE_10 0.00174526f
cc_491 N_CLKB_20 N_SE_7 0.00263447f
cc_492 N_CLKB_20 N_SE_11 0.00645061f
cc_493 N_MM1_g N_SI_5 7.546e-20
cc_494 N_CLKB_1 N_SI_5 0.000395306f
cc_495 N_CLKB_26 N_SI_5 0.000262878f
cc_496 N_CLKB_21 N_SI_7 0.000812248f
cc_497 N_CLKB_25 N_SI_6 0.000920349f
cc_498 N_CLKB_26 N_SI_6 0.00106756f
cc_499 N_CLKB_21 N_SI_5 0.00266998f
*END of SDFHx3_ASAP7_75t_R.pxi
.ENDS
** Design:	SDFHx4_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "SDFHx4_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "SDFHx4_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_SDFHx4_ASAP7_75t_R%noxref_32 VSS 1
c1 1 VSS 0.0066268f
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%NET066 VSS 2 3 1
c1 1 VSS 0.00100905f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4860 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0675 $X2=0.4860 $Y2=0.0675
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%NET067 VSS 2 3 1
c1 1 VSS 0.00101887f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0675 $X2=0.5940 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.0675 $X2=0.5940 $Y2=0.0675
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%noxref_30 VSS 1
c1 1 VSS 0.00540699f
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%noxref_31 VSS 1
c1 1 VSS 0.00554194f
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%noxref_28 VSS 1
c1 1 VSS 0.0419592f
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%noxref_29 VSS 1
c1 1 VSS 0.0419579f
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%noxref_36 VSS 1
c1 1 VSS 0.0047641f
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%noxref_40 VSS 1
c1 1 VSS 0.0423303f
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%noxref_41 VSS 1
c1 1 VSS 0.0423153f
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%noxref_38 VSS 1
c1 1 VSS 0.0417984f
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%noxref_37 VSS 1
c1 1 VSS 0.00515921f
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%noxref_39 VSS 1
c1 1 VSS 0.0418856f
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%QN VSS 31 24 25 35 36 44 45 48 49 14 16 15 13 18
+ 17 2 3 4 1
c1 1 VSS 0.0104524f
c2 2 VSS 0.0104822f
c3 3 VSS 0.00996504f
c4 4 VSS 0.00991712f
c5 13 VSS 0.00445919f
c6 14 VSS 0.00439593f
c7 15 VSS 0.00446322f
c8 16 VSS 0.00440893f
c9 17 VSS 0.019096f
c10 18 VSS 0.0200495f
c11 19 VSS 0.00795406f
c12 20 VSS 0.00328527f
c13 21 VSS 0.00333886f
r1 49 47 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.5830 $Y=0.2025 $X2=1.5805 $Y2=0.2025
r2 4 47 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.5660 $Y=0.2025 $X2=1.5805 $Y2=0.2025
r3 16 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.5515 $Y=0.2025 $X2=1.5660 $Y2=0.2025
r4 48 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.5490 $Y=0.2025 $X2=1.5515 $Y2=0.2025
r5 45 43 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.4750 $Y=0.2025 $X2=1.4725 $Y2=0.2025
r6 2 43 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.4580 $Y=0.2025 $X2=1.4725 $Y2=0.2025
r7 15 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.4435 $Y=0.2025 $X2=1.4580 $Y2=0.2025
r8 44 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.4410 $Y=0.2025 $X2=1.4435 $Y2=0.2025
r9 4 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.5660 $Y=0.2025
+ $X2=1.5660 $Y2=0.2340
r10 2 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.4580 $Y=0.2025
+ $X2=1.4580 $Y2=0.2340
r11 39 40 9.32759 $w=1.3e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=1.5660
+ $Y=0.2340 $X2=1.6060 $Y2=0.2340
r12 38 39 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.5120
+ $Y=0.2340 $X2=1.5660 $Y2=0.2340
r13 37 38 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.4580
+ $Y=0.2340 $X2=1.5120 $Y2=0.2340
r14 18 37 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=1.4480
+ $Y=0.2340 $X2=1.4580 $Y2=0.2340
r15 21 32 8.52248 $w=1.49091e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.6465 $Y=0.2340 $X2=1.6465 $Y2=0.1845
r16 21 40 7.67296 $w=1.54395e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.6465 $Y=0.2340 $X2=1.6060 $Y2=0.2340
r17 36 34 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.5830 $Y=0.0675 $X2=1.5805 $Y2=0.0675
r18 3 34 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.5660 $Y=0.0675 $X2=1.5805 $Y2=0.0675
r19 14 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.5515 $Y=0.0675 $X2=1.5660 $Y2=0.0675
r20 35 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.5490 $Y=0.0675 $X2=1.5515 $Y2=0.0675
r21 31 32 9.8736 $w=1.4e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=1.6465
+ $Y=0.1350 $X2=1.6465 $Y2=0.1845
r22 19 20 8.52248 $w=1.49091e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.6465 $Y=0.0855 $X2=1.6465 $Y2=0.0360
r23 31 19 9.8736 $w=1.4e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=1.6465
+ $Y=0.1350 $X2=1.6465 $Y2=0.0855
r24 3 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.5660 $Y=0.0675
+ $X2=1.5660 $Y2=0.0360
r25 20 30 7.67296 $w=1.54395e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.6465 $Y=0.0360 $X2=1.6060 $Y2=0.0360
r26 29 30 9.32759 $w=1.3e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=1.5660
+ $Y=0.0360 $X2=1.6060 $Y2=0.0360
r27 28 29 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.5120
+ $Y=0.0360 $X2=1.5660 $Y2=0.0360
r28 27 28 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.4580
+ $Y=0.0360 $X2=1.5120 $Y2=0.0360
r29 26 27 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=1.4480
+ $Y=0.0360 $X2=1.4580 $Y2=0.0360
r30 17 26 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.4455
+ $Y=0.0360 $X2=1.4480 $Y2=0.0360
r31 1 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.4580 $Y=0.0675
+ $X2=1.4580 $Y2=0.0360
r32 25 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.4750 $Y=0.0675 $X2=1.4725 $Y2=0.0675
r33 1 23 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.4580 $Y=0.0675 $X2=1.4725 $Y2=0.0675
r34 13 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.4435 $Y=0.0675 $X2=1.4580 $Y2=0.0675
r35 24 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.4410 $Y=0.0675 $X2=1.4435 $Y2=0.0675
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%PD3 VSS 7 9 4 5 1
c1 1 VSS 0.0103495f
c2 4 VSS 0.00189387f
c3 5 VSS 0.00311116f
r1 9 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8810 $Y=0.0675 $X2=0.8785 $Y2=0.0675
r2 5 8 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8660 $Y=0.0675 $X2=0.8785 $Y2=0.0675
r3 4 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.0675 $X2=0.8080 $Y2=0.0675
r4 7 4 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.0675 $X2=0.7955 $Y2=0.0675
r5 1 5 1e-05
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%CLK VSS 7 3 1 4 5
c1 1 VSS 0.0065664f
c2 3 VSS 0.0815892f
c3 4 VSS 0.00393737f
c4 5 VSS 0.00301133f
r1 5 8 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0720 $X2=0.0810 $Y2=0.0935
r2 7 4 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1160
r3 4 8 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1160 $X2=0.0810 $Y2=0.0935
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r5 7 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%PD4 VSS 7 9 4 5 1
c1 1 VSS 0.00859229f
c2 4 VSS 0.00181994f
c3 5 VSS 0.00311372f
r1 9 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.2050 $Y=0.2025 $X2=1.2025 $Y2=0.2025
r2 5 8 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.1900 $Y=0.2025 $X2=1.2025 $Y2=0.2025
r3 4 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.1195 $Y=0.2025 $X2=1.1320 $Y2=0.2025
r4 7 4 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.1170 $Y=0.2025 $X2=1.1195 $Y2=0.2025
r5 1 5 1e-05
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%PD5 VSS 2 4 1
c1 1 VSS 0.00096906f
r1 4 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.2050 $Y=0.0675 $X2=1.1925 $Y2=0.0675
r2 2 1 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.1710 $Y=0.0675 $X2=1.1755 $Y2=0.0675
r3 1 3 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.1755 $Y=0.0675 $X2=1.1925 $Y2=0.0675
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%MH VSS 10 39 42 50 52 13 20 18 19 4 11 15 3 17 14
+ 12 1
c1 1 VSS 0.00342262f
c2 3 VSS 0.00674529f
c3 4 VSS 0.00413327f
c4 10 VSS 0.079425f
c5 11 VSS 0.00229966f
c6 12 VSS 0.0022114f
c7 13 VSS 0.002775f
c8 14 VSS 0.000526777f
c9 15 VSS 0.000308131f
c10 16 VSS 0.000204422f
c11 17 VSS 0.0118473f
c12 18 VSS 0.00283611f
c13 19 VSS 0.000222619f
c14 20 VSS 0.000170654f
c15 21 VSS 0.00198666f
c16 22 VSS 0.00286628f
r1 52 51 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.0675 $X2=0.7705 $Y2=0.0675
r2 12 51 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7580 $Y=0.0675 $X2=0.7705 $Y2=0.0675
r3 11 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.0675 $X2=0.7000 $Y2=0.0675
r4 50 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.0675 $X2=0.6875 $Y2=0.0675
r5 3 46 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7290 $Y=0.0675
+ $X2=0.7470 $Y2=0.0900
r6 46 47 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.7470
+ $Y=0.0900 $X2=0.7470 $Y2=0.1025
r7 45 47 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.7470
+ $Y=0.1135 $X2=0.7470 $Y2=0.1025
r8 44 45 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.7470
+ $Y=0.1425 $X2=0.7470 $Y2=0.1135
r9 43 44 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.7470
+ $Y=0.1655 $X2=0.7470 $Y2=0.1425
r10 14 19 3.01468 $w=1.741e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.7470
+ $Y=0.1780 $X2=0.7470 $Y2=0.1980
r11 14 43 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.7470
+ $Y=0.1780 $X2=0.7470 $Y2=0.1655
r12 19 37 1.73214 $w=1.61034e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7470 $Y=0.1980 $X2=0.7615 $Y2=0.1980
r13 42 41 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8270 $Y=0.2025 $X2=0.8245 $Y2=0.2025
r14 40 41 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8200 $Y=0.2025 $X2=0.8245 $Y2=0.2025
r15 4 40 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8080 $Y=0.2025 $X2=0.8200 $Y2=0.2025
r16 13 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.2025 $X2=0.8080 $Y2=0.2025
r17 39 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.2025 $X2=0.7955 $Y2=0.2025
r18 36 37 1.63233 $w=1.3e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.7685
+ $Y=0.1980 $X2=0.7615 $Y2=0.1980
r19 35 36 0.816164 $w=1.3e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.7720
+ $Y=0.1980 $X2=0.7685 $Y2=0.1980
r20 34 35 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1980 $X2=0.7720 $Y2=0.1980
r21 15 20 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7965 $Y=0.1980 $X2=0.8100 $Y2=0.1980
r22 15 34 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7965
+ $Y=0.1980 $X2=0.7830 $Y2=0.1980
r23 4 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8100 $Y=0.2025
+ $X2=0.8100 $Y2=0.2160
r24 16 21 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.2160 $X2=0.8100 $Y2=0.2340
r25 16 20 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.2160 $X2=0.8100 $Y2=0.1980
r26 21 33 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.2340 $X2=0.8235 $Y2=0.2340
r27 32 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.2340 $X2=0.8235 $Y2=0.2340
r28 31 32 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.2340 $X2=0.8370 $Y2=0.2340
r29 30 31 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.2340 $X2=0.8640 $Y2=0.2340
r30 17 22 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9180 $Y=0.2340 $X2=0.9450 $Y2=0.2340
r31 17 30 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.2340 $X2=0.8910 $Y2=0.2340
r32 22 29 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.2340 $X2=0.9450 $Y2=0.2125
r33 28 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1945 $X2=0.9450 $Y2=0.2125
r34 27 28 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1780 $X2=0.9450 $Y2=0.1945
r35 26 27 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1655 $X2=0.9450 $Y2=0.1780
r36 25 26 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1540 $X2=0.9450 $Y2=0.1655
r37 24 25 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1350 $X2=0.9450 $Y2=0.1540
r38 18 24 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1160 $X2=0.9450 $Y2=0.1350
r39 10 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.9450
+ $Y=0.1350 $X2=0.9450 $Y2=0.1350
r40 1 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.9450 $Y=0.1350
+ $X2=0.9450 $Y2=0.1350
r41 3 12 1e-05
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%PD2 VSS 2 4 1
c1 1 VSS 0.000960869f
r1 4 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8810 $Y=0.2025 $X2=0.8685 $Y2=0.2025
r2 2 1 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.2025 $X2=0.8515 $Y2=0.2025
r3 1 3 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8515 $Y=0.2025 $X2=0.8685 $Y2=0.2025
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.00462576f
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%noxref_35 VSS 1
c1 1 VSS 0.0101092f
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%noxref_26 VSS 1
c1 1 VSS 0.0054357f
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.00467218f
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%noxref_27 VSS 1
c1 1 VSS 0.00546906f
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%PD1 VSS 11 21 24 8 2 9 7 1
c1 1 VSS 0.00608028f
c2 2 VSS 0.00530104f
c3 7 VSS 0.00363251f
c4 8 VSS 0.00259981f
c5 9 VSS 0.0222829f
r1 24 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.0675 $X2=0.6625 $Y2=0.0675
r2 22 23 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6580 $Y=0.0675 $X2=0.6625 $Y2=0.0675
r3 2 22 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6460 $Y=0.0675 $X2=0.6580 $Y2=0.0675
r4 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0675 $X2=0.6460 $Y2=0.0675
r5 21 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.0675 $X2=0.6335 $Y2=0.0675
r6 2 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.0675
+ $X2=0.6480 $Y2=0.0360
r7 17 18 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6255
+ $Y=0.0360 $X2=0.6480 $Y2=0.0360
r8 16 17 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6055
+ $Y=0.0360 $X2=0.6255 $Y2=0.0360
r9 15 16 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5785
+ $Y=0.0360 $X2=0.6055 $Y2=0.0360
r10 14 15 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.0360 $X2=0.5785 $Y2=0.0360
r11 13 14 13.6416 $w=1.3e-08 $l=5.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4815
+ $Y=0.0360 $X2=0.5400 $Y2=0.0360
r12 12 13 11.5429 $w=1.3e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4815 $Y2=0.0360
r13 9 12 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4205
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r14 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4320 $Y2=0.0360
r15 11 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r16 7 10 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4340 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r17 1 7 1e-05
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%noxref_34 VSS 1
c1 1 VSS 0.0108998f
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%SS VSS 9 28 32 1 12 10 11 3 14 4 17 16 13 15
c1 1 VSS 0.00417719f
c2 3 VSS 0.00854636f
c3 4 VSS 0.0063667f
c4 9 VSS 0.0814214f
c5 10 VSS 0.00423456f
c6 11 VSS 0.0046321f
c7 12 VSS 0.00145869f
c8 13 VSS 0.0019071f
c9 14 VSS 0.0010711f
c10 15 VSS 0.000441651f
c11 16 VSS 0.000684529f
c12 17 VSS 0.000442962f
r1 10 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.2815 $Y=0.0675 $X2=1.2940 $Y2=0.0675
r2 32 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.2790 $Y=0.0675 $X2=1.2815 $Y2=0.0675
r3 3 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.3055 $Y=0.0675
+ $X2=1.2960 $Y2=0.0900
r4 29 30 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.2960
+ $Y=0.0900 $X2=1.3095 $Y2=0.0900
r5 16 26 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.0900 $X2=1.3230 $Y2=0.1125
r6 16 30 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3230 $Y=0.0900 $X2=1.3095 $Y2=0.0900
r7 11 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.2815 $Y=0.2025 $X2=1.2940 $Y2=0.2025
r8 28 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.2790 $Y=0.2025 $X2=1.2815 $Y2=0.2025
r9 25 26 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.1350 $X2=1.3230 $Y2=0.1125
r10 14 17 4.8802 $w=1.615e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.1630 $X2=1.3230 $Y2=0.1910
r11 14 25 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.1630 $X2=1.3230 $Y2=0.1350
r12 4 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.2960 $Y=0.2025
+ $X2=1.2960 $Y2=0.1910
r13 17 24 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3230 $Y=0.1910 $X2=1.3095 $Y2=0.1910
r14 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.2960
+ $Y=0.1910 $X2=1.3095 $Y2=0.1910
r15 22 23 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.2850
+ $Y=0.1910 $X2=1.2960 $Y2=0.1910
r16 21 22 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.2625
+ $Y=0.1910 $X2=1.2850 $Y2=0.1910
r17 13 15 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.2330
+ $Y=0.1910 $X2=1.2150 $Y2=0.1910
r18 13 21 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=1.2330
+ $Y=0.1910 $X2=1.2625 $Y2=0.1910
r19 15 20 4.8802 $w=1.615e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.2150
+ $Y=0.1910 $X2=1.2150 $Y2=0.1630
r20 12 20 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.2150
+ $Y=0.1350 $X2=1.2150 $Y2=0.1630
r21 9 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=1.2150
+ $Y=0.1350 $X2=1.2150 $Y2=0.1350
r22 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.2150 $Y=0.1350
+ $X2=1.2150 $Y2=0.1350
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%MS VSS 11 35 39 41 43 15 1 4 17 5 3 16 13 12 14
c1 1 VSS 0.00411215f
c2 3 VSS 0.000123516f
c3 4 VSS 0.0163436f
c4 5 VSS 0.0101165f
c5 11 VSS 0.0803631f
c6 12 VSS 0.00337716f
c7 13 VSS 0.00219026f
c8 14 VSS 0.00336112f
c9 15 VSS 0.00216883f
c10 16 VSS 0.00137584f
c11 17 VSS 0.00379444f
c12 18 VSS 0.00125177f
r1 43 42 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0430 $Y=0.2025 $X2=1.0405 $Y2=0.2025
r2 15 42 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0280 $Y=0.2025 $X2=1.0405 $Y2=0.2025
r3 14 5 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9575 $Y=0.2025 $X2=0.9700 $Y2=0.2025
r4 41 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9550 $Y=0.2025 $X2=0.9575 $Y2=0.2025
r5 5 37 5.26888 $w=6.87567e-08 $l=4.85026e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9990 $Y=0.2025 $X2=0.9985 $Y2=0.1540
r6 39 38 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.0970 $Y=0.0675 $X2=1.0945 $Y2=0.0675
r7 13 38 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.0820 $Y=0.0675 $X2=1.0945 $Y2=0.0675
r8 36 37 3.71245 $w=4.12e-08 $l=1.9e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9985 $Y=0.1350 $X2=0.9985 $Y2=0.1540
r9 3 28 3.08411 $w=6.89849e-08 $l=4.86647e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9985 $Y=0.1160 $X2=1.0025 $Y2=0.0675
r10 3 36 3.71245 $w=4.12e-08 $l=1.9e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9985 $Y=0.1160 $X2=0.9985 $Y2=0.1350
r11 12 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9575 $Y=0.0675 $X2=0.9700 $Y2=0.0675
r12 35 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9550 $Y=0.0675 $X2=0.9575 $Y2=0.0675
r13 32 13 1.22083 $w=7.72e-08 $l=1.4e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.0660 $Y=0.0675 $X2=1.0800 $Y2=0.0675
r14 31 32 1.13362 $w=7.72e-08 $l=1.3e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.0530 $Y=0.0675 $X2=1.0660 $Y2=0.0675
r15 30 31 1.13362 $w=7.72e-08 $l=1.3e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.0400 $Y=0.0675 $X2=1.0530 $Y2=0.0675
r16 29 30 0.915619 $w=7.72e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.0295 $Y=0.0675 $X2=1.0400 $Y2=0.0675
r17 28 29 2.26219 $w=7.98037e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.0025 $Y=0.0675 $X2=1.0295 $Y2=0.0675
r18 27 28 1.84983 $w=8.1e-08 $l=2.25e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9800 $Y=0.0675 $X2=1.0025 $Y2=0.0675
r19 4 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.9680 $Y=0.0675
+ $X2=0.9720 $Y2=0.0720
r20 4 27 1.02647 $w=7.84667e-08 $l=1.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9680 $Y=0.0675 $X2=0.9800 $Y2=0.0675
r21 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.9585
+ $Y=0.0720 $X2=0.9720 $Y2=0.0720
r22 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.0720 $X2=0.9585 $Y2=0.0720
r23 17 18 4.75866 $w=1.41702e-08 $l=2.72259e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9180 $Y=0.0720 $X2=0.8910 $Y2=0.0755
r24 17 24 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.0720 $X2=0.9450 $Y2=0.0720
r25 18 22 3.47612 $w=1.45278e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8910 $Y=0.0755 $X2=0.8910 $Y2=0.0935
r26 16 20 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1160 $X2=0.8910 $Y2=0.1350
r27 16 22 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1160 $X2=0.8910 $Y2=0.0935
r28 11 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.8910
+ $Y=0.1350 $X2=0.8910 $Y2=0.1350
r29 1 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8910 $Y=0.1350
+ $X2=0.8910 $Y2=0.1350
r30 5 15 1e-05
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%noxref_33 VSS 1
c1 1 VSS 0.00654157f
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%D VSS 12 3 4 7 1 10 8 9 5 6
c1 1 VSS 0.00472808f
c2 3 VSS 0.0449414f
c3 4 VSS 0.00229493f
c4 5 VSS 0.00217585f
c5 6 VSS 0.00823989f
c6 7 VSS 0.00175723f
c7 8 VSS 0.00150485f
c8 9 VSS 0.00388618f
c9 10 VSS 0.00151836f
r1 6 9 3.59766 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4095
+ $Y=0.2340 $X2=0.3870 $Y2=0.2340
r2 9 17 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3870
+ $Y=0.2340 $X2=0.3870 $Y2=0.2160
r3 16 17 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3870
+ $Y=0.1980 $X2=0.3870 $Y2=0.2160
r4 15 16 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3870
+ $Y=0.1765 $X2=0.3870 $Y2=0.1980
r5 4 8 5.92955 $w=1.57138e-08 $l=3.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3870 $Y=0.1405 $X2=0.3870 $Y2=0.1080
r6 4 15 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.3870
+ $Y=0.1405 $X2=0.3870 $Y2=0.1765
r7 8 14 3.59766 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3870
+ $Y=0.1080 $X2=0.4095 $Y2=0.1080
r8 5 10 3.59766 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4365
+ $Y=0.1080 $X2=0.4590 $Y2=0.1080
r9 5 14 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4365
+ $Y=0.1080 $X2=0.4095 $Y2=0.1080
r10 12 7 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1215
r11 7 10 1.49895 $w=1.95333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1215 $X2=0.4590 $Y2=0.1080
r12 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r13 12 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1350
+ $X2=0.4590 $Y2=0.1350
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%CLKN VSS 17 18 19 20 21 93 95 12 11 28 34 1 25 27
+ 23 24 36 26 22 30 29 2 32 5 31 3 4 33 35
c1 1 VSS 0.00371175f
c2 2 VSS 8.33193e-20
c3 3 VSS 0.000297266f
c4 4 VSS 5.74436e-20
c5 5 VSS 0.000244688f
c6 11 VSS 0.00874244f
c7 12 VSS 0.00876084f
c8 17 VSS 0.0801486f
c9 18 VSS 0.00516279f
c10 19 VSS 0.00533818f
c11 20 VSS 0.00465749f
c12 21 VSS 0.0053323f
c13 22 VSS 0.00871244f
c14 23 VSS 0.00873126f
c15 24 VSS 0.00659265f
c16 25 VSS 0.0044563f
c17 26 VSS 0.00649621f
c18 27 VSS 0.0046389f
c19 28 VSS 0.00246858f
c20 29 VSS 0.000344964f
c21 30 VSS 0.00164321f
c22 31 VSS 0.00125939f
c23 32 VSS 0.0015554f
c24 33 VSS 0.0039128f
c25 34 VSS 0.00202771f
c26 35 VSS 0.0042695f
c27 36 VSS 0.0453515f
r1 95 94 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r2 23 94 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r3 93 92 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r4 22 92 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r5 12 90 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0550 $Y2=0.2340
r6 11 85 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0550 $Y2=0.0360
r7 89 90 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.2340 $X2=0.0550 $Y2=0.2340
r8 27 89 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0460 $Y2=0.2340
r9 27 35 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0180 $Y2=0.2340
r10 84 85 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.0360 $X2=0.0550 $Y2=0.0360
r11 26 84 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0460 $Y2=0.0360
r12 26 33 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0180 $Y2=0.0360
r13 35 82 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.2340 $X2=0.0180 $Y2=0.2125
r14 33 81 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0360 $X2=0.0180 $Y2=0.0540
r15 18 76 2.79569 $w=1.27128e-07 $l=5e-10 $layer=LIG $thickness=5.21026e-08
+ $X=0.6750 $Y=0.1350 $X2=0.6745 $Y2=0.1350
r16 1 73 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1440
r17 17 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r18 25 34 5.19594 $w=1.44151e-08 $l=2.80401e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1810 $X2=0.0165 $Y2=0.1530
r19 25 82 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1810 $X2=0.0180 $Y2=0.2125
r20 80 81 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0720 $X2=0.0180 $Y2=0.0540
r21 24 34 8.11081 $w=1.39615e-08 $l=4.05278e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1125 $X2=0.0165 $Y2=0.1530
r22 24 80 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1125 $X2=0.0180 $Y2=0.0720
r23 4 67 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.0530 $Y=0.1350
+ $X2=1.0530 $Y2=0.1440
r24 20 4 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=1.0530
+ $Y=0.1350 $X2=1.0530 $Y2=0.1350
r25 3 64 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8370 $Y=0.1350
+ $X2=0.8370 $Y2=0.1440
r26 19 3 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.8370
+ $Y=0.1350 $X2=0.8370 $Y2=0.1350
r27 76 77 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.6745
+ $Y=0.1350 $X2=0.6845 $Y2=0.1350
r28 2 77 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.6875 $Y=0.1350 $X2=0.6845 $Y2=0.1350
r29 2 79 5.02115 $w=1.53e-08 $l=8.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.6875
+ $Y=0.1350 $X2=0.6960 $Y2=0.1350
r30 28 73 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1160 $X2=0.1350 $Y2=0.1440
r31 70 71 1.90199 $w=1.38333e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.0255 $Y=0.1530 $X2=0.0345 $Y2=0.1530
r32 34 70 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0165
+ $Y=0.1530 $X2=0.0255 $Y2=0.1530
r33 31 67 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1160 $X2=1.0530 $Y2=0.1440
r34 30 64 10.7267 $w=1.3e-08 $l=4.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.0980 $X2=0.8370 $Y2=0.1440
r35 60 79 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6930 $Y=0.1440
+ $X2=0.6960 $Y2=0.1350
r36 29 60 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1250 $X2=0.6930 $Y2=0.1440
r37 58 59 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1530 $X2=0.1595 $Y2=0.1530
r38 58 73 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1350 $Y=0.1530
+ $X2=0.1350 $Y2=0.1440
r39 57 58 11.8927 $w=1.3e-08 $l=5.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.0840
+ $Y=0.1530 $X2=0.1350 $Y2=0.1530
r40 56 57 11.8927 $w=1.3e-08 $l=5.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.0330
+ $Y=0.1530 $X2=0.0840 $Y2=0.1530
r41 56 71 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.0330 $Y=0.1530
+ $X2=0.0345 $Y2=0.1530
r42 53 54 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M2 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1530 $X2=1.0915 $Y2=0.1530
r43 53 67 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=1.0530 $Y=0.1530
+ $X2=1.0530 $Y2=0.1440
r44 52 53 25.1845 $w=1.3e-08 $l=1.08e-07 $layer=M2 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1530 $X2=1.0530 $Y2=0.1530
r45 51 52 25.1845 $w=1.3e-08 $l=1.08e-07 $layer=M2 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1530 $X2=0.9450 $Y2=0.1530
r46 51 64 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.8370 $Y=0.1530
+ $X2=0.8370 $Y2=0.1440
r47 50 51 16.7897 $w=1.3e-08 $l=7.2e-08 $layer=M2 $thickness=3.6e-08 $X=0.7650
+ $Y=0.1530 $X2=0.8370 $Y2=0.1530
r48 49 50 16.7897 $w=1.3e-08 $l=7.2e-08 $layer=M2 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1530 $X2=0.7650 $Y2=0.1530
r49 49 60 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.6930 $Y=0.1530
+ $X2=0.6930 $Y2=0.1440
r50 48 49 61.4455 $w=1.3e-08 $l=2.635e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.4295 $Y=0.1530 $X2=0.6930 $Y2=0.1530
r51 48 59 62.9612 $w=1.3e-08 $l=2.7e-07 $layer=M2 $thickness=3.6e-08 $X=0.4295
+ $Y=0.1530 $X2=0.1595 $Y2=0.1530
r52 36 46 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=1.1365
+ $Y=0.1530 $X2=1.1610 $Y2=0.1530
r53 36 54 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M2 $thickness=3.6e-08 $X=1.1365
+ $Y=0.1530 $X2=1.0915 $Y2=0.1530
r54 43 46 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=1.1610 $Y=0.1440
+ $X2=1.1610 $Y2=0.1530
r55 32 43 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.1160 $X2=1.1610 $Y2=0.1440
r56 21 5 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=1.1610
+ $Y=0.1350 $X2=1.1610 $Y2=0.1350
r57 5 43 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.1610 $Y=0.1350
+ $X2=1.1610 $Y2=0.1440
r58 12 23 1e-05
r59 11 22 1e-05
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%PU1 VSS 12 13 24 9 2 7 1 8
c1 1 VSS 0.0047254f
c2 2 VSS 0.00474754f
c3 7 VSS 0.00221184f
c4 8 VSS 0.00219032f
c5 9 VSS 0.0164867f
r1 24 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.2025 $X2=0.7705 $Y2=0.2025
r2 8 23 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7580 $Y=0.2025 $X2=0.7705 $Y2=0.2025
r3 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7560 $Y=0.2025
+ $X2=0.7560 $Y2=0.2340
r4 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7425
+ $Y=0.2340 $X2=0.7560 $Y2=0.2340
r5 19 20 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7245
+ $Y=0.2340 $X2=0.7425 $Y2=0.2340
r6 18 19 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7065
+ $Y=0.2340 $X2=0.7245 $Y2=0.2340
r7 17 18 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.2340 $X2=0.7065 $Y2=0.2340
r8 16 17 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6730
+ $Y=0.2340 $X2=0.6930 $Y2=0.2340
r9 15 16 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.6325
+ $Y=0.2340 $X2=0.6730 $Y2=0.2340
r10 14 15 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.2340 $X2=0.6325 $Y2=0.2340
r11 9 14 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5825
+ $Y=0.2340 $X2=0.5940 $Y2=0.2340
r12 1 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2025
+ $X2=0.5940 $Y2=0.2340
r13 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.2025 $X2=0.6085 $Y2=0.2025
r14 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.2025 $X2=0.6085 $Y2=0.2025
r15 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2025 $X2=0.5940 $Y2=0.2025
r16 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.2025 $X2=0.5795 $Y2=0.2025
r17 2 8 1e-05
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%SH VSS 11 12 13 14 15 49 52 95 98 16 18 26 5 20 6
+ 17 19 2 24 1 28 23 21 22 27 29
c1 1 VSS 0.00592917f
c2 2 VSS 0.0203037f
c3 5 VSS 0.00719652f
c4 6 VSS 0.00788997f
c5 11 VSS 0.0812403f
c6 12 VSS 0.0821596f
c7 13 VSS 0.0813799f
c8 14 VSS 0.0812976f
c9 15 VSS 0.08212f
c10 16 VSS 0.00619262f
c11 17 VSS 0.00583214f
c12 18 VSS 0.0298633f
c13 19 VSS 0.0143849f
c14 20 VSS 0.00343189f
c15 21 VSS 0.011086f
c16 22 VSS 0.00429577f
c17 23 VSS 0.00429749f
c18 24 VSS 0.00321523f
c19 25 VSS 0.00358891f
c20 26 VSS 0.00167665f
c21 27 VSS 0.00505225f
c22 28 VSS 0.00146067f
c23 29 VSS 0.00478285f
r1 98 97 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0970 $Y=0.2025 $X2=1.0945 $Y2=0.2025
r2 5 97 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0820 $Y=0.2025 $X2=1.0945 $Y2=0.2025
r3 94 5 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0700 $Y=0.2025 $X2=1.0820 $Y2=0.2025
r4 17 94 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0655 $Y=0.2025 $X2=1.0700 $Y2=0.2025
r5 95 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0630 $Y=0.2025 $X2=1.0655 $Y2=0.2025
r6 5 87 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0800 $Y=0.2025
+ $X2=1.0800 $Y2=0.2340
r7 15 79 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=1.5930
+ $Y=0.1350 $X2=1.5930 $Y2=0.1350
r8 14 73 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=1.5390
+ $Y=0.1350 $X2=1.5390 $Y2=0.1350
r9 13 67 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=1.4850
+ $Y=0.1350 $X2=1.4850 $Y2=0.1350
r10 12 59 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=1.4310 $Y=0.1350 $X2=1.4310 $Y2=0.1350
r11 87 88 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.0800
+ $Y=0.2340 $X2=1.0935 $Y2=0.2340
r12 85 88 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.2340 $X2=1.0935 $Y2=0.2340
r13 84 85 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.1340
+ $Y=0.2340 $X2=1.1070 $Y2=0.2340
r14 83 84 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.2340 $X2=1.1340 $Y2=0.2340
r15 82 83 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.1880
+ $Y=0.2340 $X2=1.1610 $Y2=0.2340
r16 81 82 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.2690
+ $Y=0.2340 $X2=1.1880 $Y2=0.2340
r17 18 29 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3500 $Y=0.2340 $X2=1.3770 $Y2=0.2340
r18 18 81 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.3500
+ $Y=0.2340 $X2=1.2690 $Y2=0.2340
r19 77 79 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.5805 $Y=0.1350 $X2=1.5930 $Y2=0.1350
r20 76 77 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.5660 $Y=0.1350 $X2=1.5805 $Y2=0.1350
r21 74 76 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.5515 $Y=0.1350 $X2=1.5660 $Y2=0.1350
r22 73 74 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.5390 $Y=0.1350 $X2=1.5515 $Y2=0.1350
r23 71 73 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.5265 $Y=0.1350 $X2=1.5390 $Y2=0.1350
r24 70 71 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.5120 $Y=0.1350 $X2=1.5265 $Y2=0.1350
r25 68 70 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.4975 $Y=0.1350 $X2=1.5120 $Y2=0.1350
r26 67 68 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.4850 $Y=0.1350 $X2=1.4975 $Y2=0.1350
r27 65 67 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.4725 $Y=0.1350 $X2=1.4850 $Y2=0.1350
r28 64 65 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.4580 $Y=0.1350 $X2=1.4725 $Y2=0.1350
r29 62 64 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.4435 $Y=0.1350 $X2=1.4580 $Y2=0.1350
r30 60 62 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=1.4405 $Y=0.1350 $X2=1.4435 $Y2=0.1350
r31 59 60 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=1.4310
+ $Y=0.1350 $X2=1.4405 $Y2=0.1350
r32 2 59 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=1.4215
+ $Y=0.1350 $X2=1.4310 $Y2=0.1350
r33 29 55 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3770 $Y=0.2340 $X2=1.3770 $Y2=0.2125
r34 56 59 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.4310 $Y=0.1350
+ $X2=1.4310 $Y2=0.1350
r35 24 56 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.4040
+ $Y=0.1350 $X2=1.4310 $Y2=0.1350
r36 24 28 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.4040 $Y=0.1350 $X2=1.3770 $Y2=0.1350
r37 23 28 7.44771 $w=1.42162e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3770 $Y=0.1720 $X2=1.3770 $Y2=0.1350
r38 23 55 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=1.3770
+ $Y=0.1720 $X2=1.3770 $Y2=0.2125
r39 28 54 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.3770
+ $Y=0.1350 $X2=1.3770 $Y2=0.1125
r40 53 54 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.3770
+ $Y=0.0900 $X2=1.3770 $Y2=0.1125
r41 22 27 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3770 $Y=0.0630 $X2=1.3770 $Y2=0.0360
r42 22 53 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.3770
+ $Y=0.0630 $X2=1.3770 $Y2=0.0900
r43 52 51 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.1510 $Y=0.0675 $X2=1.1485 $Y2=0.0675
r44 50 51 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.1440 $Y=0.0675 $X2=1.1485 $Y2=0.0675
r45 6 50 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.1320 $Y=0.0675 $X2=1.1440 $Y2=0.0675
r46 16 6 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.1195 $Y=0.0675 $X2=1.1320 $Y2=0.0675
r47 49 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.1170 $Y=0.0675 $X2=1.1195 $Y2=0.0675
r48 27 47 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3770 $Y=0.0360 $X2=1.3500 $Y2=0.0360
r49 6 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.1340 $Y=0.0675
+ $X2=1.1340 $Y2=0.0360
r50 46 47 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=1.3095
+ $Y=0.0360 $X2=1.3500 $Y2=0.0360
r51 45 46 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=1.2850
+ $Y=0.0360 $X2=1.3095 $Y2=0.0360
r52 21 25 3.60008 $w=1.51951e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.2715 $Y=0.0360 $X2=1.2510 $Y2=0.0360
r53 21 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.2715
+ $Y=0.0360 $X2=1.2850 $Y2=0.0360
r54 42 43 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.1340
+ $Y=0.0360 $X2=1.1475 $Y2=0.0360
r55 40 43 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0360 $X2=1.1475 $Y2=0.0360
r56 39 40 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.1880
+ $Y=0.0360 $X2=1.1610 $Y2=0.0360
r57 38 39 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.2150
+ $Y=0.0360 $X2=1.1880 $Y2=0.0360
r58 19 25 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.2330
+ $Y=0.0360 $X2=1.2510 $Y2=0.0360
r59 19 38 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.2330
+ $Y=0.0360 $X2=1.2150 $Y2=0.0360
r60 25 37 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.2510
+ $Y=0.0360 $X2=1.2510 $Y2=0.0540
r61 36 37 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.2510
+ $Y=0.0665 $X2=1.2510 $Y2=0.0540
r62 35 36 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.2510
+ $Y=0.0755 $X2=1.2510 $Y2=0.0665
r63 34 35 3.38125 $w=1.3e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=1.2510
+ $Y=0.0900 $X2=1.2510 $Y2=0.0755
r64 33 34 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.2510
+ $Y=0.1025 $X2=1.2510 $Y2=0.0900
r65 20 26 3.2503 $w=1.53684e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.2510 $Y=0.1160 $X2=1.2510 $Y2=0.1350
r66 20 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.2510
+ $Y=0.1160 $X2=1.2510 $Y2=0.1025
r67 26 31 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.2510
+ $Y=0.1350 $X2=1.2690 $Y2=0.1350
r68 11 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=1.2690
+ $Y=0.1350 $X2=1.2690 $Y2=0.1350
r69 1 31 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.2690 $Y=0.1350
+ $X2=1.2690 $Y2=0.1350
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%SI VSS 14 3 12 9 1 4 8 7 5 10 6
c1 1 VSS 0.00311798f
c2 3 VSS 0.0068723f
c3 4 VSS 0.00154003f
c4 5 VSS 0.00159569f
c5 6 VSS 0.00171696f
c6 7 VSS 0.00176022f
c7 8 VSS 0.00716307f
c8 9 VSS 0.00167574f
c9 10 VSS 0.00162732f
c10 11 VSS 0.003537f
c11 12 VSS 0.00158821f
r1 8 11 3.59766 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.7245
+ $Y=0.0360 $X2=0.7020 $Y2=0.0360
r2 7 12 2.45586 $w=1.44e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.0540 $X2=0.7020 $Y2=0.0665
r3 7 11 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.0540 $X2=0.7020 $Y2=0.0360
r4 12 19 1.40651 $w=1.51875e-08 $l=1.45774e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7020 $Y=0.0665 $X2=0.6885 $Y2=0.0720
r5 18 19 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.6730
+ $Y=0.0720 $X2=0.6885 $Y2=0.0720
r6 6 10 1.03257 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6595 $Y=0.0720 $X2=0.6480 $Y2=0.0720
r7 6 18 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6595
+ $Y=0.0720 $X2=0.6730 $Y2=0.0720
r8 5 17 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6480 $Y=0.0935 $X2=0.6480 $Y2=0.1150
r9 5 10 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6480 $Y=0.0935 $X2=0.6480 $Y2=0.0720
r10 16 17 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6345 $Y=0.1150 $X2=0.6480 $Y2=0.1150
r11 9 16 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.1150 $X2=0.6345 $Y2=0.1150
r12 14 4 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1250
r13 4 9 1.15159 $w=1.75e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1250 $X2=0.6210 $Y2=0.1150
r14 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1350
r15 14 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6210 $Y=0.1350
+ $X2=0.6210 $Y2=0.1350
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%NET54 VSS 15 34 35 37 12 3 13 11 2 10 1
c1 1 VSS 0.00606074f
c2 2 VSS 0.00604706f
c3 3 VSS 0.0034366f
c4 10 VSS 0.00447676f
c5 11 VSS 0.00333157f
c6 12 VSS 0.00265957f
c7 13 VSS 0.00532717f
r1 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.2025 $X2=0.6460 $Y2=0.2025
r2 37 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.2025 $X2=0.6335 $Y2=0.2025
r3 35 33 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r4 2 33 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5400 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r5 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.2025 $X2=0.5400 $Y2=0.2025
r6 34 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.2025 $X2=0.5255 $Y2=0.2025
r7 3 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.2025
+ $X2=0.6480 $Y2=0.1980
r8 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.2025
+ $X2=0.5400 $Y2=0.1980
r9 29 30 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6345
+ $Y=0.1980 $X2=0.6480 $Y2=0.1980
r10 28 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1980 $X2=0.6345 $Y2=0.1980
r11 27 28 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.6055
+ $Y=0.1980 $X2=0.6210 $Y2=0.1980
r12 26 27 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.5895
+ $Y=0.1980 $X2=0.6055 $Y2=0.1980
r13 25 26 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5780
+ $Y=0.1980 $X2=0.5895 $Y2=0.1980
r14 24 25 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1980 $X2=0.5780 $Y2=0.1980
r15 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5535
+ $Y=0.1980 $X2=0.5670 $Y2=0.1980
r16 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1980 $X2=0.5535 $Y2=0.1980
r17 21 22 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5265
+ $Y=0.1980 $X2=0.5400 $Y2=0.1980
r18 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1980 $X2=0.5265 $Y2=0.1980
r19 19 20 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.1980 $X2=0.5130 $Y2=0.1980
r20 18 19 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4635
+ $Y=0.1980 $X2=0.4860 $Y2=0.1980
r21 17 18 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4545
+ $Y=0.1980 $X2=0.4635 $Y2=0.1980
r22 16 17 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4455
+ $Y=0.1980 $X2=0.4545 $Y2=0.1980
r23 13 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.1980 $X2=0.4455 $Y2=0.1980
r24 1 13 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.1980
r25 15 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r26 10 14 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4340 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r27 1 10 1e-05
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%SE VSS 24 5 6 8 14 7 12 13 9 15 10 11 1 2
c1 1 VSS 0.0104652f
c2 2 VSS 0.00464909f
c3 5 VSS 0.0823582f
c4 6 VSS 0.0450049f
c5 7 VSS 0.00521658f
c6 8 VSS 0.00390567f
c7 9 VSS 0.00181048f
c8 10 VSS 0.00368449f
c9 11 VSS 0.00669263f
c10 12 VSS 0.00159082f
c11 13 VSS 0.00747562f
c12 14 VSS 0.00224836f
c13 15 VSS 0.00718839f
r1 2 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1350
+ $X2=0.5670 $Y2=0.1350
r2 6 2 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1350
r3 14 30 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.5670 $Y=0.0720 $X2=0.5670
+ $Y2=0.0810
r4 35 36 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1250 $X2=0.5670 $Y2=0.1350
r5 34 35 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1150 $X2=0.5670 $Y2=0.1250
r6 33 34 3.96423 $w=1.3e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0980 $X2=0.5670 $Y2=0.1150
r7 10 33 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0855 $X2=0.5670 $Y2=0.0980
r8 10 30 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.5670 $Y=0.0855 $X2=0.5670
+ $Y2=0.0810
r9 10 14 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.0855 $X2=0.5670 $Y2=0.0720
r10 29 30 37.7767 $w=1.3e-08 $l=1.62e-07 $layer=M2 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0810 $X2=0.5670 $Y2=0.0810
r11 28 29 37.7767 $w=1.3e-08 $l=1.62e-07 $layer=M2 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0810 $X2=0.4050 $Y2=0.0810
r12 15 28 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.2315
+ $Y=0.0810 $X2=0.2430 $Y2=0.0810
r13 8 12 10.3626 $w=1.39091e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.1845 $X2=0.2430 $Y2=0.1350
r14 8 13 10.3626 $w=1.39091e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.1845 $X2=0.2430 $Y2=0.2340
r15 25 26 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0810 $X2=0.2430 $Y2=0.1080
r16 25 28 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.2430 $Y=0.0810
+ $X2=0.2430 $Y2=0.0810
r17 7 25 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0585 $X2=0.2430 $Y2=0.0810
r18 7 11 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0585 $X2=0.2430 $Y2=0.0360
r19 12 26 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2430 $Y2=0.1080
r20 24 9 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2800
+ $Y=0.1350 $X2=0.2615 $Y2=0.1350
r21 9 12 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2615 $Y=0.1350 $X2=0.2430 $Y2=0.1350
r22 24 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2800 $Y=0.1350
+ $X2=0.2765 $Y2=0.1350
r23 20 22 4.72579 $w=1.53e-08 $l=8e-09 $layer=LIG $thickness=4.8e-08 $X=0.2845
+ $Y=0.1350 $X2=0.2765 $Y2=0.1350
r24 1 19 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.2880
+ $Y=0.1350 $X2=0.2980 $Y2=0.1350
r25 1 20 1.73797 $w=1.72143e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.2880 $Y=0.1350 $X2=0.2845 $Y2=0.1350
r26 5 19 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2980 $Y2=0.1350
r27 5 20 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2845 $Y2=0.1350
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%CLKB VSS 11 12 55 57 5 19 21 16 6 15 1 18 2 14 13
+ 17 20
c1 1 VSS 0.000156357f
c2 2 VSS 0.000133017f
c3 5 VSS 0.00772697f
c4 6 VSS 0.00852242f
c5 11 VSS 0.00433513f
c6 12 VSS 0.00444025f
c7 13 VSS 0.00910614f
c8 14 VSS 0.00916086f
c9 15 VSS 0.00577509f
c10 16 VSS 0.00333338f
c11 17 VSS 0.000812397f
c12 18 VSS 0.00176199f
c13 19 VSS 0.0064026f
c14 20 VSS 0.00248124f
c15 21 VSS 0.0293127f
r1 13 5 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0675 $X2=0.1600 $Y2=0.0675
r2 57 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1475 $Y2=0.0675
r3 14 6 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1600 $Y2=0.2025
r4 55 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r5 5 50 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0675
+ $X2=0.1620 $Y2=0.0360
r6 6 47 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r7 50 51 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r8 15 50 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1505
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r9 47 48 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r10 19 45 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2340 $X2=0.1890 $Y2=0.2125
r11 19 48 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2340 $X2=0.1755 $Y2=0.2340
r12 20 41 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.1890 $Y2=0.0540
r13 20 51 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1755 $Y2=0.0360
r14 1 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7830 $Y=0.1350
+ $X2=0.7830 $Y2=0.1260
r15 11 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.7830
+ $Y=0.1350 $X2=0.7830 $Y2=0.1350
r16 44 45 11.5429 $w=1.3e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1630 $X2=0.1890 $Y2=0.2125
r17 43 44 10.7267 $w=1.3e-08 $l=4.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1170 $X2=0.1890 $Y2=0.1630
r18 42 43 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1070 $X2=0.1890 $Y2=0.1170
r19 40 41 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0720 $X2=0.1890 $Y2=0.0540
r20 16 40 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0935 $X2=0.1890 $Y2=0.0720
r21 16 42 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0935 $X2=0.1890 $Y2=0.1070
r22 17 38 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.0890 $X2=0.7830 $Y2=0.1260
r23 36 37 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1170 $X2=0.2135 $Y2=0.1170
r24 36 43 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1890 $Y=0.1170
+ $X2=0.1890 $Y2=0.1170
r25 34 37 44.6558 $w=1.3e-08 $l=1.915e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.4050 $Y=0.1170 $X2=0.2135 $Y2=0.1170
r26 31 32 37.7767 $w=1.3e-08 $l=1.62e-07 $layer=M2 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1170 $X2=1.1070 $Y2=0.1170
r27 30 31 37.7767 $w=1.3e-08 $l=1.62e-07 $layer=M2 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1170 $X2=0.9450 $Y2=0.1170
r28 30 38 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.7830 $Y=0.1170
+ $X2=0.7830 $Y2=0.1260
r29 21 30 24.6015 $w=1.3e-08 $l=1.055e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.6775 $Y=0.1170 $X2=0.7830 $Y2=0.1170
r30 21 34 63.5442 $w=1.3e-08 $l=2.725e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.6775 $Y=0.1170 $X2=0.4050 $Y2=0.1170
r31 26 32 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=1.1070 $Y=0.1260
+ $X2=1.1070 $Y2=0.1170
r32 18 26 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.1070 $X2=1.1070 $Y2=0.1260
r33 12 2 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=1.1070
+ $Y=0.1350 $X2=1.1070 $Y2=0.1350
r34 2 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.1070 $Y=0.1350
+ $X2=1.1070 $Y2=0.1260
.ends

.subckt PM_SDFHx4_ASAP7_75t_R%SEN VSS 9 37 39 10 16 17 11 4 1 19 3 13 15 14
c1 1 VSS 0.00392879f
c2 3 VSS 0.00773156f
c3 4 VSS 0.00804802f
c4 9 VSS 0.081547f
c5 10 VSS 0.0052735f
c6 11 VSS 0.00529801f
c7 12 VSS 0.000481334f
c8 13 VSS 0.00263259f
c9 14 VSS 0.00346815f
c10 15 VSS 0.00286126f
c11 16 VSS 0.00688966f
c12 17 VSS 0.00655501f
c13 18 VSS 0.000260545f
c14 19 VSS 0.000605237f
r1 11 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3220 $Y2=0.2025
r2 39 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r3 10 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3220 $Y2=0.0675
r4 37 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r5 4 34 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.2340
r6 3 31 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0675
+ $X2=0.3240 $Y2=0.0360
r7 34 35 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.2340 $X2=0.3375 $Y2=0.2340
r8 17 29 10.3626 $w=1.39091e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.2340 $X2=0.3510 $Y2=0.1845
r9 17 35 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.2340 $X2=0.3375 $Y2=0.2340
r10 31 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.0360 $X2=0.3375 $Y2=0.0360
r11 16 32 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.0360 $X2=0.3375 $Y2=0.0360
r12 28 29 11.5429 $w=1.3e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1845
r13 27 28 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1125 $X2=0.3510 $Y2=0.1350
r14 13 18 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0900 $X2=0.3510 $Y2=0.0720
r15 13 27 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0900 $X2=0.3510 $Y2=0.1125
r16 12 18 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0540 $X2=0.3510 $Y2=0.0720
r17 12 16 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0540 $X2=0.3510 $Y2=0.0360
r18 18 26 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0720 $X2=0.3690 $Y2=0.0720
r19 25 26 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.3980
+ $Y=0.0720 $X2=0.3690 $Y2=0.0720
r20 24 25 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4430
+ $Y=0.0720 $X2=0.3980 $Y2=0.0720
r21 14 19 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4860 $Y=0.0720 $X2=0.5130 $Y2=0.0720
r22 14 24 10.0272 $w=1.3e-08 $l=4.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.0720 $X2=0.4430 $Y2=0.0720
r23 19 23 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0720 $X2=0.5130 $Y2=0.0900
r24 15 21 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1125 $X2=0.5130 $Y2=0.1350
r25 15 23 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1125 $X2=0.5130 $Y2=0.0900
r26 9 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r27 1 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.1350
+ $X2=0.5130 $Y2=0.1350
.ends


*
.SUBCKT SDFHx4_ASAP7_75t_R VSS VDD CLK SE D SI QN
*
* VSS VSS
* VDD VDD
* CLK CLK
* SE SE
* D D
* SI SI
* QN QN
*
*

MM20 N_MM20_d N_MM20_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM23 N_MM23_d N_MM23_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM30 N_MM30_d N_MM31_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM29 N_MM29_d N_MM26_g N_MM29_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM28 N_MM28_d N_MM0_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM27 N_MM27_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM2_g N_MM5_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM1_g N_MM9_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM6_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM12 N_MM12_d N_MM12_g N_MM12_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM17 N_MM17_d N_MM17_g N_MM17_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM16 N_MM16_d N_MM16_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM14 N_MM14_d N_MM14_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24 N_MM24_d N_MM24_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@4 N_MM24@4_d N_MM24@4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@3 N_MM24@3_d N_MM24@3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@2 N_MM24@2_d N_MM24@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM21 N_MM21_d N_MM20_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM22 N_MM22_d N_MM23_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM31 N_MM31_d N_MM31_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM26 N_MM26_d N_MM26_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g N_MM3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g N_MM2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM6_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM13 N_MM13_d N_MM13_g N_MM13_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM18 N_MM18_d N_MM12_g N_MM18_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM19 N_MM19_d N_MM16_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM15 N_MM15_d N_MM14_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25 N_MM25_d N_MM24_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@4 N_MM25@4_d N_MM24@4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@3 N_MM25@3_d N_MM24@3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@2 N_MM25@2_d N_MM24@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "SDFHx4_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "SDFHx4_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_SDFHx4_ASAP7_75t_R%noxref_32 VSS N_noxref_32_1
+ PM_SDFHx4_ASAP7_75t_R%noxref_32
cc_1 N_noxref_32_1 N_MM26_g 0.00151698f
cc_2 N_noxref_32_1 N_SEN_10 0.000920687f
cc_3 N_noxref_32_1 N_PD1_7 0.0354609f
cc_4 N_noxref_32_1 N_noxref_30_1 0.00766401f
x_PM_SDFHx4_ASAP7_75t_R%NET066 VSS N_MM29_s N_MM28_d N_NET066_1
+ PM_SDFHx4_ASAP7_75t_R%NET066
cc_5 N_NET066_1 N_MM26_g 0.0172883f
cc_6 N_NET066_1 N_MM0_g 0.0172804f
x_PM_SDFHx4_ASAP7_75t_R%NET067 VSS N_MM27_d N_MM5_s N_NET067_1
+ PM_SDFHx4_ASAP7_75t_R%NET067
cc_7 N_NET067_1 N_MM3_g 0.0173966f
cc_8 N_NET067_1 N_MM2_g 0.0172783f
x_PM_SDFHx4_ASAP7_75t_R%noxref_30 VSS N_noxref_30_1
+ PM_SDFHx4_ASAP7_75t_R%noxref_30
cc_9 N_noxref_30_1 N_MM31_g 0.00134085f
cc_10 N_noxref_30_1 N_SEN_10 0.0378036f
x_PM_SDFHx4_ASAP7_75t_R%noxref_31 VSS N_noxref_31_1
+ PM_SDFHx4_ASAP7_75t_R%noxref_31
cc_11 N_noxref_31_1 N_MM31_g 0.00134383f
cc_12 N_noxref_31_1 N_SEN_11 0.0376784f
cc_13 N_noxref_31_1 N_noxref_30_1 0.00122999f
x_PM_SDFHx4_ASAP7_75t_R%noxref_28 VSS N_noxref_28_1
+ PM_SDFHx4_ASAP7_75t_R%noxref_28
cc_14 N_noxref_28_1 N_MM31_g 0.00180328f
cc_15 N_noxref_28_1 N_CLKB_5 0.000133462f
cc_16 N_noxref_28_1 N_CLKB_13 0.000671416f
cc_17 N_noxref_28_1 N_noxref_26_1 0.00765072f
x_PM_SDFHx4_ASAP7_75t_R%noxref_29 VSS N_noxref_29_1
+ PM_SDFHx4_ASAP7_75t_R%noxref_29
cc_18 N_noxref_29_1 N_MM31_g 0.00179844f
cc_19 N_noxref_29_1 N_CLKB_6 0.000135924f
cc_20 N_noxref_29_1 N_CLKB_14 0.000674258f
cc_21 N_noxref_29_1 N_noxref_27_1 0.00765311f
cc_22 N_noxref_29_1 N_noxref_28_1 0.00122493f
x_PM_SDFHx4_ASAP7_75t_R%noxref_36 VSS N_noxref_36_1
+ PM_SDFHx4_ASAP7_75t_R%noxref_36
cc_23 N_noxref_36_1 N_SS_3 0.00145621f
cc_24 N_noxref_36_1 N_SS_10 0.0374735f
cc_25 N_noxref_36_1 N_MM14_g 0.00152626f
x_PM_SDFHx4_ASAP7_75t_R%noxref_40 VSS N_noxref_40_1
+ PM_SDFHx4_ASAP7_75t_R%noxref_40
cc_26 N_noxref_40_1 N_MM24@2_g 0.00147423f
cc_27 N_noxref_40_1 N_QN_14 0.000832699f
x_PM_SDFHx4_ASAP7_75t_R%noxref_41 VSS N_noxref_41_1
+ PM_SDFHx4_ASAP7_75t_R%noxref_41
cc_28 N_noxref_41_1 N_MM24@2_g 0.00146661f
cc_29 N_noxref_41_1 N_QN_16 0.000832498f
cc_30 N_noxref_41_1 N_noxref_40_1 0.00177139f
x_PM_SDFHx4_ASAP7_75t_R%noxref_38 VSS N_noxref_38_1
+ PM_SDFHx4_ASAP7_75t_R%noxref_38
cc_31 N_noxref_38_1 N_SS_10 0.00110149f
cc_32 N_noxref_38_1 N_MM24_g 0.00176105f
cc_33 N_noxref_38_1 N_noxref_36_1 0.00753653f
x_PM_SDFHx4_ASAP7_75t_R%noxref_37 VSS N_noxref_37_1
+ PM_SDFHx4_ASAP7_75t_R%noxref_37
cc_34 N_noxref_37_1 N_SS_11 0.0377243f
cc_35 N_noxref_37_1 N_MM14_g 0.00168082f
cc_36 N_noxref_37_1 N_noxref_36_1 0.00121773f
x_PM_SDFHx4_ASAP7_75t_R%noxref_39 VSS N_noxref_39_1
+ PM_SDFHx4_ASAP7_75t_R%noxref_39
cc_37 N_noxref_39_1 N_SS_11 0.000808725f
cc_38 N_noxref_39_1 N_MM24_g 0.00180988f
cc_39 N_noxref_39_1 N_noxref_37_1 0.00766121f
cc_40 N_noxref_39_1 N_noxref_38_1 0.00124117f
x_PM_SDFHx4_ASAP7_75t_R%QN VSS QN N_MM24_d N_MM24@4_d N_MM24@3_d N_MM24@2_d
+ N_MM25_d N_MM25@4_d N_MM25@3_d N_MM25@2_d N_QN_14 N_QN_16 N_QN_15 N_QN_13
+ N_QN_18 N_QN_17 N_QN_2 N_QN_3 N_QN_4 N_QN_1 PM_SDFHx4_ASAP7_75t_R%QN
cc_41 N_QN_14 N_SH_27 0.000154126f
cc_42 N_QN_14 N_SH_29 0.00016251f
cc_43 N_QN_14 N_MM24_g 0.000360622f
cc_44 N_QN_14 N_SH_22 0.000443736f
cc_45 N_QN_14 N_SH_23 0.000470506f
cc_46 N_QN_14 N_SH_2 0.00123424f
cc_47 N_QN_16 N_MM24@3_g 0.0305524f
cc_48 N_QN_15 N_MM24_g 0.0305192f
cc_49 N_QN_13 N_MM24_g 0.067239f
cc_50 N_QN_18 N_MM24@3_g 0.00090569f
cc_51 N_QN_17 N_MM24@3_g 0.000940779f
cc_52 N_QN_2 N_SH_24 0.00100245f
cc_53 N_QN_3 N_MM24@3_g 0.00176823f
cc_54 N_QN_4 N_MM24@3_g 0.00182077f
cc_55 N_QN_1 N_MM24_g 0.00208974f
cc_56 N_QN_2 N_MM24_g 0.00213295f
cc_57 N_QN_15 N_SH_2 0.00972117f
cc_58 N_QN_14 N_MM24@2_g 0.0367225f
cc_59 N_QN_13 N_MM24@4_g 0.0367759f
cc_60 N_QN_14 N_MM24@3_g 0.0676825f
x_PM_SDFHx4_ASAP7_75t_R%PD3 VSS N_MM9_s N_MM8_d N_PD3_4 N_PD3_5 N_PD3_1
+ PM_SDFHx4_ASAP7_75t_R%PD3
cc_61 N_PD3_4 N_CLKN_3 0.00189226f
cc_62 N_PD3_4 N_CLKN_30 0.001064f
cc_63 N_PD3_4 N_MM10_g 0.0740883f
cc_64 N_PD3_4 N_CLKB_17 0.000525719f
cc_65 N_PD3_4 N_CLKB_1 0.000623541f
cc_66 N_PD3_4 N_MM1_g 0.03465f
cc_67 N_PD3_5 N_MM11_g 0.0366661f
cc_68 N_PD3_1 N_MH_3 0.00120033f
cc_69 N_PD3_1 N_MH_12 0.00288579f
x_PM_SDFHx4_ASAP7_75t_R%CLK VSS CLK N_MM20_g N_CLK_1 N_CLK_4 N_CLK_5
+ PM_SDFHx4_ASAP7_75t_R%CLK
x_PM_SDFHx4_ASAP7_75t_R%PD4 VSS N_MM18_s N_MM19_d N_PD4_4 N_PD4_5 N_PD4_1
+ PM_SDFHx4_ASAP7_75t_R%PD4
cc_70 N_PD4_4 N_CLKN_31 5.85084e-20
cc_71 N_PD4_4 N_CLKN_5 0.00225618f
cc_72 N_PD4_4 N_CLKN_32 0.000995784f
cc_73 N_PD4_4 N_MM17_g 0.073678f
cc_74 N_PD4_4 N_CLKB_18 0.000203209f
cc_75 N_PD4_4 N_CLKB_2 0.000694531f
cc_76 N_PD4_4 N_MM12_g 0.0342011f
cc_77 N_PD4_5 N_SS_1 0.000812342f
cc_78 N_PD4_5 N_MM16_g 0.0351091f
cc_79 N_PD4_1 N_SH_5 0.00135725f
cc_80 N_PD4_1 N_SH_17 0.00115519f
cc_81 N_PD4_1 N_SH_18 0.00447388f
x_PM_SDFHx4_ASAP7_75t_R%PD5 VSS N_MM17_s N_MM16_d N_PD5_1
+ PM_SDFHx4_ASAP7_75t_R%PD5
cc_82 N_PD5_1 N_MM17_g 0.0170138f
cc_83 N_PD5_1 N_MM16_g 0.0170874f
x_PM_SDFHx4_ASAP7_75t_R%MH VSS N_MM6_g N_MM1_d N_MM10_d N_MM4_d N_MM9_d N_MH_13
+ N_MH_20 N_MH_18 N_MH_19 N_MH_4 N_MH_11 N_MH_15 N_MH_3 N_MH_17 N_MH_14 N_MH_12
+ N_MH_1 PM_SDFHx4_ASAP7_75t_R%MH
cc_84 N_MH_13 N_CLKN_31 4.13386e-20
cc_85 N_MH_13 N_MM13_g 4.40212e-20
cc_86 N_MH_13 N_CLKN_4 4.43965e-20
cc_87 N_MH_13 N_CLKN_36 0.000224847f
cc_88 N_MH_13 N_CLKN_30 0.000342541f
cc_89 N_MH_13 N_CLKN_29 0.000302321f
cc_90 N_MH_20 N_CLKN_30 0.000924849f
cc_91 N_MH_18 N_CLKN_31 0.000287308f
cc_92 N_MH_19 N_CLKN_29 0.000310655f
cc_93 N_MH_4 N_CLKN_3 0.000339259f
cc_94 N_MH_11 N_MM4_g 0.0346616f
cc_95 N_MH_15 N_CLKN_30 0.000464687f
cc_96 N_MH_3 N_CLKN_2 0.000832119f
cc_97 N_MH_13 N_CLKN_3 0.00085154f
cc_98 N_MH_17 N_CLKN_30 0.000892325f
cc_99 N_MH_14 N_CLKN_36 0.000928093f
cc_100 N_MH_4 N_CLKN_30 0.0010206f
cc_101 N_MH_4 N_MM10_g 0.00125079f
cc_102 N_MH_3 N_MM4_g 0.00172392f
cc_103 N_MH_11 N_CLKN_2 0.00197899f
cc_104 N_MH_14 N_CLKN_29 0.00310036f
cc_105 N_MH_18 N_CLKN_36 0.00344676f
cc_106 N_MH_13 N_MM10_g 0.0351614f
cc_107 N_MH_14 N_SI_7 0.000383051f
cc_108 N_MH_14 N_SI_8 0.00149895f
cc_109 N_MH_3 N_SI_12 0.00179191f
cc_110 N_MH_14 N_SI_12 0.00334305f
cc_111 N_MH_12 N_CLKB_17 0.000975678f
cc_112 N_MH_13 N_MM1_g 0.0155852f
cc_113 N_MH_15 N_CLKB_17 0.000759234f
cc_114 N_MH_4 N_MM1_g 0.000896563f
cc_115 N_MH_14 N_CLKB_1 0.00096818f
cc_116 N_MH_3 N_MM1_g 0.00117981f
cc_117 N_MH_13 N_CLKB_1 0.00161434f
cc_118 N_MH_18 N_CLKB_21 0.00207726f
cc_119 N_MH_14 N_CLKB_17 0.00872816f
cc_120 N_MH_12 N_MM1_g 0.053549f
cc_121 N_MH_1 N_MS_12 0.000472131f
cc_122 N_MH_1 N_MS_1 0.000583955f
cc_123 N_MM6_g N_MS_4 0.000913329f
cc_124 N_MH_18 N_MS_17 0.000982872f
cc_125 N_MH_1 N_MS_3 0.00261736f
cc_126 N_MM6_g N_MS_5 0.0017653f
cc_127 N_MM6_g N_MM11_g 0.00188084f
cc_128 N_MH_1 N_MS_14 0.00219472f
cc_129 N_MM6_g N_MS_14 0.0147562f
cc_130 N_MH_18 N_MS_16 0.00535186f
cc_131 N_MM6_g N_MS_12 0.0560734f
x_PM_SDFHx4_ASAP7_75t_R%PD2 VSS N_MM10_s N_MM11_d N_PD2_1
+ PM_SDFHx4_ASAP7_75t_R%PD2
cc_132 N_PD2_1 N_MM10_g 0.0170064f
cc_133 N_PD2_1 N_MM11_g 0.017083f
x_PM_SDFHx4_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_SDFHx4_ASAP7_75t_R%noxref_25
cc_134 N_noxref_25_1 N_MM20_g 0.00145212f
cc_135 N_noxref_25_1 N_CLKN_22 0.000131175f
cc_136 N_noxref_25_1 N_CLKN_35 5.74907e-20
cc_137 N_noxref_25_1 N_CLKN_34 6.85133e-20
cc_138 N_noxref_25_1 N_CLKN_11 7.53042e-20
cc_139 N_noxref_25_1 N_CLKN_24 0.000125616f
cc_140 N_noxref_25_1 N_CLKN_25 0.000179511f
cc_141 N_noxref_25_1 N_CLKN_12 0.00049868f
cc_142 N_noxref_25_1 N_CLKN_23 0.0373367f
cc_143 N_noxref_25_1 N_noxref_24_1 0.00175969f
x_PM_SDFHx4_ASAP7_75t_R%noxref_35 VSS N_noxref_35_1
+ PM_SDFHx4_ASAP7_75t_R%noxref_35
cc_144 N_noxref_35_1 N_MM13_g 0.0100763f
cc_145 N_noxref_35_1 N_MS_5 0.000890787f
cc_146 N_noxref_35_1 N_MS_3 0.0014053f
cc_147 N_noxref_35_1 N_MS_4 0.00210579f
cc_148 N_noxref_35_1 N_MS_12 0.016313f
cc_149 N_noxref_35_1 N_MS_15 0.0163095f
cc_150 N_noxref_35_1 N_MS_14 0.0781059f
cc_151 N_noxref_35_1 N_MM6_g 0.00325707f
x_PM_SDFHx4_ASAP7_75t_R%noxref_26 VSS N_noxref_26_1
+ PM_SDFHx4_ASAP7_75t_R%noxref_26
cc_152 N_noxref_26_1 N_MM23_g 0.00135812f
cc_153 N_noxref_26_1 N_CLKB_16 0.000112077f
cc_154 N_noxref_26_1 N_CLKB_5 0.000418458f
cc_155 N_noxref_26_1 N_CLKB_13 0.0372249f
x_PM_SDFHx4_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_SDFHx4_ASAP7_75t_R%noxref_24
cc_156 N_noxref_24_1 N_MM20_g 0.00145517f
cc_157 N_noxref_24_1 N_CLKN_23 0.000133675f
cc_158 N_noxref_24_1 N_CLKN_34 4.64767e-20
cc_159 N_noxref_24_1 N_CLKN_25 5.52438e-20
cc_160 N_noxref_24_1 N_CLKN_33 5.62629e-20
cc_161 N_noxref_24_1 N_CLKN_12 7.35668e-20
cc_162 N_noxref_24_1 N_CLKN_24 0.000263193f
cc_163 N_noxref_24_1 N_CLKN_11 0.000505587f
cc_164 N_noxref_24_1 N_CLKN_22 0.0373987f
x_PM_SDFHx4_ASAP7_75t_R%noxref_27 VSS N_noxref_27_1
+ PM_SDFHx4_ASAP7_75t_R%noxref_27
cc_165 N_noxref_27_1 N_MM23_g 0.00136017f
cc_166 N_noxref_27_1 N_CLKB_16 0.000110919f
cc_167 N_noxref_27_1 N_CLKB_6 0.000413219f
cc_168 N_noxref_27_1 N_CLKB_14 0.0371717f
cc_169 N_noxref_27_1 N_noxref_26_1 0.0012378f
x_PM_SDFHx4_ASAP7_75t_R%PD1 VSS N_MM29_d N_MM5_d N_MM4_s N_PD1_8 N_PD1_2
+ N_PD1_9 N_PD1_7 N_PD1_1 PM_SDFHx4_ASAP7_75t_R%PD1
cc_170 N_PD1_8 N_CLKN_2 0.000826798f
cc_171 N_PD1_8 N_CLKN_36 0.000135212f
cc_172 N_PD1_2 N_MM4_g 0.000776244f
cc_173 N_PD1_8 N_MM4_g 0.0333589f
cc_174 N_PD1_9 N_SE_10 0.000494535f
cc_175 N_PD1_9 N_MM3_g 0.00023683f
cc_176 N_PD1_9 N_SE_15 0.000899365f
cc_177 N_PD1_9 N_SE_14 0.00599414f
cc_178 N_PD1_7 N_D_1 0.000790732f
cc_179 N_PD1_1 N_MM26_g 0.00172411f
cc_180 N_PD1_7 N_MM26_g 0.0351919f
cc_181 N_PD1_9 N_MM0_g 0.000241587f
cc_182 N_PD1_1 N_SEN_14 0.00183166f
cc_183 N_PD1_9 N_SEN_14 0.00454406f
cc_184 N_PD1_9 N_SEN_19 0.00666503f
cc_185 N_PD1_8 N_SI_5 0.000348966f
cc_186 N_PD1_2 N_SI_10 0.000382294f
cc_187 N_PD1_8 N_SI_1 0.000670386f
cc_188 N_PD1_9 N_SI_6 0.000750406f
cc_189 N_PD1_9 N_SI_10 0.00119559f
cc_190 N_PD1_9 N_SI_9 0.00188155f
cc_191 N_PD1_2 N_MM2_g 0.00195849f
cc_192 N_PD1_8 N_MM2_g 0.035085f
cc_193 N_PD1_8 N_MH_11 0.000556245f
cc_194 N_PD1_2 N_MH_3 0.00116368f
cc_195 N_PD1_8 N_MH_3 0.00216711f
x_PM_SDFHx4_ASAP7_75t_R%noxref_34 VSS N_noxref_34_1
+ PM_SDFHx4_ASAP7_75t_R%noxref_34
cc_196 N_noxref_34_1 N_MM4_g 0.00507028f
cc_197 N_noxref_34_1 N_CLKN_2 0.00678357f
cc_198 N_noxref_34_1 N_MM1_g 0.00347983f
cc_199 N_noxref_34_1 N_MH_3 0.00112779f
cc_200 N_noxref_34_1 N_MH_12 0.0166195f
cc_201 N_noxref_34_1 N_MH_11 0.0563743f
cc_202 N_noxref_34_1 N_PU1_8 0.0368508f
x_PM_SDFHx4_ASAP7_75t_R%SS VSS N_MM16_g N_MM15_d N_MM14_d N_SS_1 N_SS_12
+ N_SS_10 N_SS_11 N_SS_3 N_SS_14 N_SS_4 N_SS_17 N_SS_16 N_SS_13 N_SS_15
+ PM_SDFHx4_ASAP7_75t_R%SS
cc_203 N_MM16_g N_CLKN_32 0.000766597f
cc_204 N_MM16_g N_CLKN_36 0.000409187f
cc_205 N_SS_1 N_CLKN_5 0.00230703f
cc_206 N_SS_12 N_CLKN_32 0.00322945f
cc_207 N_MM16_g N_MM17_g 0.00512898f
x_PM_SDFHx4_ASAP7_75t_R%MS VSS N_MM11_g N_MM6_d N_MM12_d N_MM7_d N_MM13_d
+ N_MS_15 N_MS_1 N_MS_4 N_MS_17 N_MS_5 N_MS_3 N_MS_16 N_MS_13 N_MS_12 N_MS_14
+ PM_SDFHx4_ASAP7_75t_R%MS
cc_208 N_MS_15 N_MM17_g 5.14858e-20
cc_209 N_MS_15 N_CLKN_31 0.000113613f
cc_210 N_MS_15 N_CLKN_30 0.000570366f
cc_211 N_MS_1 N_CLKN_3 0.00213434f
cc_212 N_MS_4 N_CLKN_4 0.00404991f
cc_213 N_MS_17 N_CLKN_36 0.00116281f
cc_214 N_MS_5 N_MM13_g 0.00146895f
cc_215 N_MS_3 N_CLKN_4 0.00149343f
cc_216 N_MS_5 N_CLKN_31 0.0016739f
cc_217 N_MS_16 N_CLKN_30 0.00363601f
cc_218 N_MS_4 N_MM13_g 0.00460967f
cc_219 N_MM11_g N_MM10_g 0.00494641f
cc_220 N_MS_13 N_MM13_g 0.0166959f
cc_221 N_MS_15 N_MM13_g 0.0557837f
cc_222 N_MS_13 N_MM1_g 5.8916e-20
cc_223 N_MS_13 N_CLKB_2 0.000917397f
cc_224 N_MS_13 N_CLKB_21 0.000229421f
cc_225 N_MS_13 N_CLKB_18 0.000699016f
cc_226 N_MS_17 N_CLKB_21 0.00076153f
cc_227 N_MS_4 N_MM12_g 0.0015885f
cc_228 N_MS_16 N_CLKB_21 0.00246682f
cc_229 N_MS_13 N_MM12_g 0.0344599f
x_PM_SDFHx4_ASAP7_75t_R%noxref_33 VSS N_noxref_33_1
+ PM_SDFHx4_ASAP7_75t_R%noxref_33
cc_230 N_noxref_33_1 N_MM26_g 0.00165339f
cc_231 N_noxref_33_1 N_SEN_11 0.000814771f
cc_232 N_noxref_33_1 N_NET54_10 0.0355325f
cc_233 N_noxref_33_1 N_noxref_31_1 0.0076476f
cc_234 N_noxref_33_1 N_noxref_32_1 0.00123858f
x_PM_SDFHx4_ASAP7_75t_R%D VSS D N_MM26_g N_D_4 N_D_7 N_D_1 N_D_10 N_D_8 N_D_9
+ N_D_5 N_D_6 PM_SDFHx4_ASAP7_75t_R%D
cc_235 N_D_4 N_CLKN_36 0.00150305f
cc_236 N_D_7 N_CLKN_36 0.00213543f
x_PM_SDFHx4_ASAP7_75t_R%CLKN VSS N_MM23_g N_MM4_g N_MM10_g N_MM13_g N_MM17_g
+ N_MM20_d N_MM21_d N_CLKN_12 N_CLKN_11 N_CLKN_28 N_CLKN_34 N_CLKN_1 N_CLKN_25
+ N_CLKN_27 N_CLKN_23 N_CLKN_24 N_CLKN_36 N_CLKN_26 N_CLKN_22 N_CLKN_30
+ N_CLKN_29 N_CLKN_2 N_CLKN_32 N_CLKN_5 N_CLKN_31 N_CLKN_3 N_CLKN_4 N_CLKN_33
+ N_CLKN_35 PM_SDFHx4_ASAP7_75t_R%CLKN
cc_237 N_CLKN_12 N_MM20_g 0.00146129f
cc_238 N_CLKN_11 N_MM20_g 0.00162425f
cc_239 N_CLKN_28 N_MM20_g 0.000218069f
cc_240 N_CLKN_34 N_MM20_g 0.000260444f
cc_241 N_CLKN_1 N_MM20_g 0.000384055f
cc_242 N_CLKN_25 N_MM20_g 0.000404132f
cc_243 N_CLKN_27 N_MM20_g 0.000435529f
cc_244 N_CLKN_23 N_MM20_g 0.0156443f
cc_245 N_CLKN_1 N_CLK_1 0.000471728f
cc_246 N_CLKN_24 N_CLK_4 0.000983719f
cc_247 N_CLKN_36 N_CLK_4 0.00113949f
cc_248 N_CLKN_12 N_CLK_1 0.00118881f
cc_249 N_MM23_g N_MM20_g 0.00164698f
cc_250 N_CLKN_28 N_CLK_4 0.00192333f
cc_251 N_CLKN_23 N_CLK_1 0.00200473f
cc_252 N_CLKN_26 N_CLK_5 0.00403559f
cc_253 N_CLKN_34 N_CLK_4 0.00763457f
cc_254 N_CLKN_22 N_MM20_g 0.0554627f
x_PM_SDFHx4_ASAP7_75t_R%PU1 VSS N_MM3_d N_MM2_d N_MM1_s N_PU1_9 N_PU1_2 N_PU1_7
+ N_PU1_1 N_PU1_8 PM_SDFHx4_ASAP7_75t_R%PU1
cc_255 N_PU1_9 N_MM10_g 7.60872e-20
cc_256 N_PU1_9 N_CLKN_2 0.000406134f
cc_257 N_PU1_9 N_MM4_g 0.000496161f
cc_258 N_PU1_2 N_MM4_g 0.000472533f
cc_259 N_PU1_9 N_CLKN_36 0.000618699f
cc_260 N_PU1_9 N_CLKN_29 0.00154168f
cc_261 N_PU1_7 N_SE_2 0.000657751f
cc_262 N_PU1_1 N_MM3_g 0.00091539f
cc_263 N_PU1_7 N_MM3_g 0.0338741f
cc_264 N_PU1_7 N_SI_1 0.000667918f
cc_265 N_PU1_1 N_MM2_g 0.000914446f
cc_266 N_PU1_7 N_MM2_g 0.0338744f
cc_267 N_PU1_8 N_CLKB_21 0.000192735f
cc_268 N_PU1_8 N_CLKB_1 0.000958692f
cc_269 N_PU1_2 N_MM1_g 0.000919812f
cc_270 N_PU1_8 N_MM1_g 0.0337223f
cc_271 N_PU1_8 N_MH_13 0.00124889f
cc_272 N_PU1_2 N_MH_14 0.000703887f
cc_273 N_PU1_2 N_MH_15 0.000729373f
cc_274 N_PU1_9 N_MH_15 0.0011781f
cc_275 N_PU1_2 N_MH_4 0.00353749f
cc_276 N_PU1_9 N_MH_19 0.00467199f
cc_277 N_PU1_7 N_NET54_13 0.000559739f
cc_278 N_PU1_7 N_NET54_12 0.000639861f
cc_279 N_PU1_1 N_NET54_13 0.000664062f
cc_280 N_PU1_7 N_NET54_11 0.00112618f
cc_281 N_PU1_1 N_NET54_3 0.00185531f
cc_282 N_PU1_1 N_NET54_2 0.00429339f
cc_283 N_PU1_9 N_NET54_13 0.00985101f
x_PM_SDFHx4_ASAP7_75t_R%SH VSS N_MM14_g N_MM24_g N_MM24@4_g N_MM24@3_g
+ N_MM24@2_g N_MM12_s N_MM17_d N_MM13_s N_MM18_d N_SH_16 N_SH_18 N_SH_26 N_SH_5
+ N_SH_20 N_SH_6 N_SH_17 N_SH_19 N_SH_2 N_SH_24 N_SH_1 N_SH_28 N_SH_23 N_SH_21
+ N_SH_22 N_SH_27 N_SH_29 PM_SDFHx4_ASAP7_75t_R%SH
cc_284 N_SH_16 N_CLKN_32 8.31206e-20
cc_285 N_SH_16 N_CLKN_31 6.52414e-20
cc_286 N_SH_18 N_CLKN_32 0.00282826f
cc_287 N_SH_26 N_CLKN_32 0.000160244f
cc_288 N_SH_5 N_CLKN_31 0.00155812f
cc_289 N_SH_20 N_CLKN_32 0.000207034f
cc_290 N_SH_5 N_CLKN_4 0.000222946f
cc_291 N_SH_6 N_CLKN_5 0.000332798f
cc_292 N_SH_17 N_MM13_g 0.0345578f
cc_293 N_SH_19 N_CLKN_32 0.000615262f
cc_294 N_SH_17 N_CLKN_4 0.000717349f
cc_295 N_SH_16 N_CLKN_5 0.000862353f
cc_296 N_SH_18 N_CLKN_36 0.0010089f
cc_297 N_SH_5 N_MM13_g 0.00132631f
cc_298 N_SH_6 N_MM17_g 0.00137626f
cc_299 N_SH_6 N_CLKN_32 0.00193937f
cc_300 N_SH_16 N_MM17_g 0.0353999f
cc_301 N_SH_16 N_CLKB_18 8.80643e-20
cc_302 N_SH_6 N_CLKB_18 0.00197109f
cc_303 N_SH_18 N_CLKB_18 0.000330453f
cc_304 N_SH_18 N_CLKB_21 0.00039058f
cc_305 N_SH_17 N_MM12_g 0.0155755f
cc_306 N_SH_5 N_CLKB_2 0.000423625f
cc_307 N_SH_5 N_MM12_g 0.000981121f
cc_308 N_SH_19 N_CLKB_18 0.0010272f
cc_309 N_SH_6 N_MM12_g 0.00128879f
cc_310 N_SH_17 N_CLKB_2 0.00135155f
cc_311 N_SH_16 N_MM12_g 0.05378f
cc_312 N_SH_18 N_MS_4 0.000171735f
cc_313 N_SH_5 N_MS_4 0.00017938f
cc_314 N_SH_19 N_MS_4 0.000192698f
cc_315 N_SH_6 N_MS_4 0.00141622f
cc_316 N_SH_17 N_MS_4 0.000568709f
cc_317 N_SH_17 N_MS_15 0.000612187f
cc_318 N_SH_16 N_MS_13 0.000613524f
cc_319 N_SH_5 N_MS_5 0.00125521f
cc_320 N_SH_17 N_MS_5 0.00149883f
cc_321 N_SH_16 N_MS_4 0.00240463f
cc_322 N_SH_16 N_SS_10 9.15269e-20
cc_323 N_SH_2 N_SS_10 9.54403e-20
cc_324 N_SH_24 N_SS_10 0.000152189f
cc_325 N_SH_6 N_SS_10 0.000228342f
cc_326 N_SH_18 N_SS_10 0.000440877f
cc_327 N_SH_19 N_SS_10 0.000442266f
cc_328 N_MM14_g N_SS_11 0.0158137f
cc_329 N_SH_1 N_SS_1 0.000591203f
cc_330 N_SH_26 N_SS_1 0.000631315f
cc_331 N_SH_20 N_SS_3 0.000695555f
cc_332 N_SH_28 N_SS_14 0.000743323f
cc_333 N_SH_1 N_SS_4 0.0012544f
cc_334 N_SH_18 N_SS_17 0.00140842f
cc_335 N_SH_23 N_SS_17 0.00143701f
cc_336 N_MM14_g N_SS_4 0.00170784f
cc_337 N_MM14_g N_MM16_g 0.00192283f
cc_338 N_SH_21 N_SS_16 0.00201129f
cc_339 N_SH_1 N_SS_11 0.00215211f
cc_340 N_MM14_g N_SS_3 0.00244116f
cc_341 N_SH_22 N_SS_16 0.00248973f
cc_342 N_SH_20 N_SS_12 0.00272761f
cc_343 N_SH_26 N_SS_14 0.00319257f
cc_344 N_SH_26 N_SS_16 0.00325462f
cc_345 N_SH_18 N_SS_13 0.00329539f
cc_346 N_SH_26 N_SS_12 0.00426691f
cc_347 N_SH_18 N_SS_15 0.00556963f
cc_348 N_MM14_g N_SS_10 0.0557687f
x_PM_SDFHx4_ASAP7_75t_R%SI VSS SI N_MM2_g N_SI_12 N_SI_9 N_SI_1 N_SI_4 N_SI_8
+ N_SI_7 N_SI_5 N_SI_10 N_SI_6 PM_SDFHx4_ASAP7_75t_R%SI
cc_349 N_MM2_g N_CLKN_30 6.44155e-20
cc_350 N_MM2_g N_CLKN_36 8.36984e-20
cc_351 N_MM2_g N_CLKN_29 0.000733614f
cc_352 N_MM2_g N_CLKN_2 0.000207368f
cc_353 N_SI_12 N_CLKN_29 0.000300056f
cc_354 N_SI_9 N_CLKN_2 0.000310765f
cc_355 N_SI_1 N_CLKN_2 0.000966796f
cc_356 N_SI_4 N_CLKN_36 0.0014133f
cc_357 N_SI_9 N_CLKN_29 0.00180084f
cc_358 N_MM2_g N_MM4_g 0.00343911f
cc_359 N_MM2_g N_SE_14 0.000232133f
cc_360 N_SI_4 N_SE_10 0.000608625f
cc_361 N_SI_1 N_SE_2 0.00210804f
cc_362 N_SI_9 N_SE_10 0.00111156f
cc_363 N_SI_9 N_SE_14 0.00152511f
cc_364 N_MM2_g N_MM3_g 0.00543653f
x_PM_SDFHx4_ASAP7_75t_R%NET54 VSS N_MM26_d N_MM0_d N_MM3_s N_MM2_s N_NET54_12
+ N_NET54_3 N_NET54_13 N_NET54_11 N_NET54_2 N_NET54_10 N_NET54_1
+ PM_SDFHx4_ASAP7_75t_R%NET54
cc_365 N_NET54_12 N_CLKN_29 0.000807935f
cc_366 N_NET54_12 N_CLKN_2 0.000999375f
cc_367 N_NET54_3 N_MM4_g 0.00117671f
cc_368 N_NET54_13 N_CLKN_36 0.0038341f
cc_369 N_NET54_12 N_MM4_g 0.0360709f
cc_370 N_NET54_11 N_SE_2 0.00102596f
cc_371 N_NET54_2 N_MM3_g 0.000840499f
cc_372 N_NET54_13 N_SE_10 0.00239954f
cc_373 N_NET54_11 N_MM3_g 0.0335087f
cc_374 N_NET54_10 N_D_6 0.00072493f
cc_375 N_NET54_10 N_D_1 0.000785024f
cc_376 N_NET54_13 N_D_4 0.00143216f
cc_377 N_NET54_1 N_MM26_g 0.00185507f
cc_378 N_NET54_13 N_D_6 0.00233081f
cc_379 N_NET54_13 N_D_7 0.00473115f
cc_380 N_NET54_10 N_MM26_g 0.0342561f
cc_381 N_NET54_11 N_SEN_1 0.000902991f
cc_382 N_NET54_2 N_MM0_g 0.000865107f
cc_383 N_NET54_13 N_SEN_15 0.0022396f
cc_384 N_NET54_11 N_MM0_g 0.0343778f
cc_385 N_NET54_12 N_SI_1 0.000706888f
cc_386 N_NET54_3 N_MM2_g 0.000918109f
cc_387 N_NET54_13 N_SI_4 0.00214602f
cc_388 N_NET54_12 N_MM2_g 0.0337008f
x_PM_SDFHx4_ASAP7_75t_R%SE VSS SE N_MM31_g N_MM3_g N_SE_8 N_SE_14 N_SE_7
+ N_SE_12 N_SE_13 N_SE_9 N_SE_15 N_SE_10 N_SE_11 N_SE_1 N_SE_2
+ PM_SDFHx4_ASAP7_75t_R%SE
cc_389 N_SE_8 N_CLKN_28 7.26176e-20
cc_390 N_SE_8 N_CLKN_26 2.09559e-20
cc_391 N_SE_8 N_CLKN_24 2.69027e-20
cc_392 N_SE_8 N_CLKN_1 4.30473e-20
cc_393 N_SE_8 N_MM4_g 5.13684e-20
cc_394 N_SE_14 N_CLKN_36 6.14828e-20
cc_395 N_SE_7 N_CLKN_36 0.000145116f
cc_396 N_SE_12 N_CLKN_36 0.000195653f
cc_397 N_SE_13 N_CLKN_36 0.000257688f
cc_398 N_SE_9 N_CLKN_36 0.000406826f
cc_399 N_SE_15 N_CLKN_36 0.00116707f
cc_400 N_SE_10 N_CLKN_36 0.00160727f
cc_401 N_SE_8 N_CLKN_36 0.00313343f
x_PM_SDFHx4_ASAP7_75t_R%CLKB VSS N_MM1_g N_MM12_g N_MM22_d N_MM23_d N_CLKB_5
+ N_CLKB_19 N_CLKB_21 N_CLKB_16 N_CLKB_6 N_CLKB_15 N_CLKB_1 N_CLKB_18 N_CLKB_2
+ N_CLKB_14 N_CLKB_13 N_CLKB_17 N_CLKB_20 PM_SDFHx4_ASAP7_75t_R%CLKB
cc_402 N_CLKB_5 N_CLK_5 0.000160779f
cc_403 N_CLKB_19 N_CLK_5 5.85481e-20
cc_404 N_CLKB_21 N_CLK_5 6.76808e-20
cc_405 N_CLKB_16 N_CLK_5 0.000162254f
cc_406 N_CLKB_6 N_CLK_5 0.000276037f
cc_407 N_CLKB_15 N_CLK_5 0.00140024f
cc_408 N_CLKB_21 N_CLKN_11 2.50275e-20
cc_409 N_CLKB_21 N_MM4_g 3.49927e-20
cc_410 N_CLKB_21 N_CLKN_28 3.81724e-20
cc_411 N_CLKB_21 N_CLKN_27 4.80315e-20
cc_412 N_CLKB_15 N_CLKN_24 5.89049e-20
cc_413 N_CLKB_1 N_CLKN_2 0.000142841f
cc_414 N_CLKB_5 N_MM23_g 0.00120133f
cc_415 N_CLKB_6 N_CLKN_28 0.000175169f
cc_416 N_CLKB_18 N_CLKN_32 0.00177579f
cc_417 N_CLKB_21 N_CLKN_29 0.000637095f
cc_418 N_CLKB_16 N_CLKN_28 0.00648893f
cc_419 N_CLKB_2 N_CLKN_5 0.000818871f
cc_420 N_CLKB_21 N_CLKN_31 0.000437184f
cc_421 N_CLKB_14 N_MM23_g 0.0157674f
cc_422 N_CLKB_13 N_MM23_g 0.0537713f
cc_423 N_CLKB_17 N_CLKN_36 0.000527447f
cc_424 N_CLKB_21 N_CLKN_30 0.000582056f
cc_425 N_CLKB_6 N_CLKN_1 0.000754531f
cc_426 N_CLKB_19 N_CLKN_28 0.000777063f
cc_427 N_CLKB_16 N_CLKN_36 0.000795625f
cc_428 N_CLKB_15 N_CLKN_26 0.000798299f
cc_429 N_CLKB_1 N_CLKN_3 0.00167085f
cc_430 N_CLKB_18 N_CLKN_36 0.000883522f
cc_431 N_CLKB_2 N_CLKN_4 0.00241793f
cc_432 N_CLKB_6 N_MM23_g 0.00135091f
cc_433 N_MM12_g N_MM17_g 0.00163458f
cc_434 N_CLKB_13 N_CLKN_1 0.00165759f
cc_435 N_MM1_g N_MM10_g 0.00333693f
cc_436 N_CLKB_17 N_CLKN_30 0.00424613f
cc_437 N_MM12_g N_MM13_g 0.00496365f
cc_438 N_CLKB_18 N_CLKN_31 0.00523573f
cc_439 N_CLKB_21 N_CLKN_36 0.0748413f
cc_440 N_CLKB_16 N_SE_15 0.00020681f
cc_441 N_CLKB_15 N_SE_15 9.74764e-20
cc_442 N_CLKB_5 N_SE_7 0.000182783f
cc_443 N_CLKB_6 N_SE_8 0.000190267f
cc_444 N_CLKB_16 N_SE_7 0.00233398f
cc_445 N_CLKB_21 N_SE_10 0.000835869f
cc_446 N_CLKB_21 N_SE_14 0.000342413f
cc_447 N_CLKB_21 N_SE_9 0.000399849f
cc_448 N_CLKB_21 N_SE_7 0.000654674f
cc_449 N_CLKB_19 N_SE_13 0.000850896f
cc_450 N_CLKB_20 N_SE_11 0.000887766f
cc_451 N_CLKB_16 N_SE_8 0.00168764f
cc_452 N_CLKB_16 N_SE_12 0.00427242f
cc_453 N_CLKB_21 N_SE_15 0.0282124f
cc_454 N_CLKB_21 N_D_5 0.00244749f
cc_455 N_CLKB_21 N_SI_12 0.000270167f
cc_456 N_CLKB_21 N_SI_8 0.000983432f
cc_457 N_CLKB_17 N_SI_8 0.00101131f
cc_458 N_CLKB_21 N_SI_9 0.00232947f
x_PM_SDFHx4_ASAP7_75t_R%SEN VSS N_MM0_g N_MM30_d N_MM31_d N_SEN_10 N_SEN_16
+ N_SEN_17 N_SEN_11 N_SEN_4 N_SEN_1 N_SEN_19 N_SEN_3 N_SEN_13 N_SEN_15 N_SEN_14
+ PM_SDFHx4_ASAP7_75t_R%SEN
cc_459 N_SEN_10 N_SE_11 0.000151975f
cc_460 N_SEN_10 N_SE_15 0.000738822f
cc_461 N_SEN_16 N_SE_7 0.000317471f
cc_462 N_SEN_17 N_SE_8 0.000337038f
cc_463 N_SEN_11 N_MM31_g 0.0157623f
cc_464 N_SEN_4 N_SE_1 0.000590479f
cc_465 N_SEN_1 N_SE_2 0.00157418f
cc_466 N_SEN_19 N_SE_14 0.000770639f
cc_467 N_SEN_17 N_SE_13 0.000808123f
cc_468 N_SEN_16 N_SE_11 0.00106618f
cc_469 N_SEN_4 N_MM31_g 0.00109792f
cc_470 N_SEN_3 N_MM31_g 0.00111958f
cc_471 N_SEN_13 N_SE_9 0.00198221f
cc_472 N_SEN_11 N_SE_1 0.00204653f
cc_473 N_SEN_15 N_SE_10 0.00305448f
cc_474 N_MM0_g N_MM3_g 0.00327844f
cc_475 N_SEN_14 N_SE_15 0.00413679f
cc_476 N_SEN_10 N_MM31_g 0.0543721f
cc_477 N_SEN_1 N_D_1 0.00220925f
cc_478 N_SEN_14 N_D_10 0.00121323f
cc_479 N_SEN_13 N_D_8 0.00134983f
cc_480 N_SEN_17 N_D_9 0.00170642f
cc_481 N_SEN_15 N_D_7 0.00191981f
cc_482 N_MM0_g N_MM26_g 0.00499343f
cc_483 N_SEN_14 N_D_5 0.00646648f
cc_484 N_SEN_13 N_D_4 0.00904751f
*END of SDFHx4_ASAP7_75t_R.pxi
.ENDS
** Design:	SDFLx1_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "SDFLx1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "SDFLx1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_SDFLx1_ASAP7_75t_R%NET0167 VSS 2 3 1
c1 1 VSS 0.000993624f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3780 $Y2=0.0675
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%NET0144 VSS 12 13 27 28 9 7 1 8 2
c1 1 VSS 0.00544179f
c2 2 VSS 0.00525369f
c3 7 VSS 0.00333871f
c4 8 VSS 0.00335752f
c5 9 VSS 0.00273131f
r1 28 26 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r2 2 26 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r4 27 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r5 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4280 $Y2=0.1980
r6 21 22 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4185
+ $Y=0.1980 $X2=0.4280 $Y2=0.1980
r7 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1980 $X2=0.4185 $Y2=0.1980
r8 19 20 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.3875
+ $Y=0.1980 $X2=0.4050 $Y2=0.1980
r9 18 19 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3695
+ $Y=0.1980 $X2=0.3875 $Y2=0.1980
r10 17 18 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1980 $X2=0.3695 $Y2=0.1980
r11 16 17 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.1980 $X2=0.3510 $Y2=0.1980
r12 15 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1980 $X2=0.3375 $Y2=0.1980
r13 14 15 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3130
+ $Y=0.1980 $X2=0.3240 $Y2=0.1980
r14 9 14 0.699569 $w=1.3e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.3100
+ $Y=0.1980 $X2=0.3130 $Y2=0.1980
r15 1 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.1980
r16 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r17 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r18 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r19 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.00418148f
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.00417137f
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%noxref_30 VSS 1
c1 1 VSS 0.0126736f
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%PD4 VSS 2 4 1
c1 1 VSS 0.0010217f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9890 $Y=0.2295 $X2=0.9765 $Y2=0.2295
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9550 $Y=0.2295 $X2=0.9595 $Y2=0.2295
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9595 $Y=0.2295 $X2=0.9765 $Y2=0.2295
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%PD3 VSS 2 4 1
c1 1 VSS 0.000909455f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.0405 $X2=0.7065 $Y2=0.0405
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.0405 $X2=0.6895 $Y2=0.0405
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6895 $Y=0.0405 $X2=0.7065 $Y2=0.0405
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%PD2 VSS 7 12 5 1 4
c1 1 VSS 0.00739927f
c2 4 VSS 0.00184482f
c3 5 VSS 0.00233019f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7040 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r3 9 5 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.6765
+ $Y=0.2295 $X2=0.7020 $Y2=0.2295
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.6615
+ $Y=0.2295 $X2=0.6765 $Y2=0.2295
r5 1 8 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.6480
+ $Y=0.2295 $X2=0.6615 $Y2=0.2295
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.2295 $X2=0.6460 $Y2=0.2295
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.2295 $X2=0.6335 $Y2=0.2295
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%CLK VSS 11 3 4 6 1 5
c1 1 VSS 0.00304854f
c2 3 VSS 0.0599119f
c3 4 VSS 0.00147271f
c4 5 VSS 0.00465386f
c5 6 VSS 0.00195426f
r1 5 14 4.60559 $w=1.39091e-08 $l=2.74591e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0630 $X2=0.1030 $Y2=0.0900
r2 13 14 1.45753 $w=1.53529e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.0900 $X2=0.1030 $Y2=0.0900
r3 6 13 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0900 $X2=0.0945 $Y2=0.0900
r4 11 10 0.757867 $w=1.3e-08 $l=3.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1500 $X2=0.0810 $Y2=0.1467
r5 9 10 2.73998 $w=1.3e-08 $l=1.17e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1467
r6 8 9 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1235 $X2=0.0810 $Y2=0.1350
r7 4 8 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1100 $X2=0.0810 $Y2=0.1235
r8 4 6 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1100 $X2=0.0810 $Y2=0.0900
r9 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r10 1 9 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%noxref_34 VSS 1
c1 1 VSS 0.00481257f
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%noxref_33 VSS 1
c1 1 VSS 0.00413925f
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%PU1 VSS 13 24 26 10 2 11 8 1 9
c1 1 VSS 0.00669234f
c2 2 VSS 0.00872161f
c3 8 VSS 0.00352464f
c4 9 VSS 0.00233431f
c5 10 VSS 0.00218811f
c6 11 VSS 0.0218062f
r1 26 25 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r2 10 25 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5420 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r3 9 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4840 $Y2=0.2025
r4 24 9 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r5 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5130 $Y=0.2025
+ $X2=0.4900 $Y2=0.2340
r6 20 21 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4810
+ $Y=0.2340 $X2=0.4900 $Y2=0.2340
r7 19 20 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4690
+ $Y=0.2340 $X2=0.4810 $Y2=0.2340
r8 18 19 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4540
+ $Y=0.2340 $X2=0.4690 $Y2=0.2340
r9 17 18 17.7224 $w=1.3e-08 $l=7.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.4540 $Y2=0.2340
r10 16 17 19.5879 $w=1.3e-08 $l=8.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2940
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r11 15 16 5.59655 $w=1.3e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.2940 $Y2=0.2340
r12 11 15 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2580
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r13 8 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2160
+ $X2=0.2700 $Y2=0.2340
r14 1 8 23.8708 $w=2.02e-08 $l=4.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.2700 $Y=0.1755 $X2=0.2700 $Y2=0.2160
r15 13 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r16 8 12 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r17 2 10 1e-05
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%noxref_27 VSS 1
c1 1 VSS 0.00438459f
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%noxref_29 VSS 1
c1 1 VSS 0.00572578f
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%noxref_28 VSS 1
c1 1 VSS 0.00558406f
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%D VSS 4 3 1 5
c1 1 VSS 0.0077051f
c2 3 VSS 0.0462888f
c3 4 VSS 0.00470479f
c4 5 VSS 0.00374569f
r1 5 7 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.1080 $X2=0.4050 $Y2=0.1215
r2 4 7 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1215
r3 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r4 4 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%noxref_26 VSS 1
c1 1 VSS 0.00439643f
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%SI VSS 14 3 5 6 7 4 1
c1 1 VSS 0.00616603f
c2 3 VSS 0.00750067f
c3 4 VSS 0.00328232f
c4 5 VSS 0.00322923f
c5 6 VSS 0.00369854f
c6 7 VSS 0.00388018f
r1 6 19 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1980 $X2=0.5130 $Y2=0.1765
r2 5 7 3.2503 $w=1.53684e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1540 $X2=0.5130 $Y2=0.1350
r3 5 19 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1540 $X2=0.5130 $Y2=0.1765
r4 7 16 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1350 $X2=0.4945 $Y2=0.1350
r5 15 16 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4845
+ $Y=0.1350 $X2=0.4945 $Y2=0.1350
r6 14 15 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4750
+ $Y=0.1350 $X2=0.4845 $Y2=0.1350
r7 14 4 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4750
+ $Y=0.1350 $X2=0.4635 $Y2=0.1350
r8 14 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4750 $Y=0.1350
+ $X2=0.4790 $Y2=0.1350
r9 11 12 4.43042 $w=1.53e-08 $l=7.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.4715
+ $Y=0.1350 $X2=0.4790 $Y2=0.1350
r10 9 11 1.86855 $w=1.78125e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.4675 $Y=0.1350 $X2=0.4715 $Y2=0.1350
r11 1 9 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.4575
+ $Y=0.1350 $X2=0.4675 $Y2=0.1350
r12 3 1 2.53453 $w=1.32811e-07 $l=1.5e-09 $layer=LIG $thickness=5.23243e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4575 $Y2=0.1350
r13 3 11 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4715 $Y2=0.1350
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%NET0168 VSS 14 27 7 9 1 11 12 10 2 8
c1 1 VSS 0.00638167f
c2 2 VSS 0.0056662f
c3 7 VSS 0.004629f
c4 8 VSS 0.0031536f
c5 9 VSS 0.000879202f
c6 10 VSS 0.0174797f
c7 11 VSS 0.00124295f
c8 12 VSS 0.00198915f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0675 $X2=0.4840 $Y2=0.0675
r2 27 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4715 $Y2=0.0675
r3 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0675
+ $X2=0.4860 $Y2=0.0360
r4 23 24 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4475
+ $Y=0.0360 $X2=0.4860 $Y2=0.0360
r5 22 23 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4070
+ $Y=0.0360 $X2=0.4475 $Y2=0.0360
r6 21 22 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.3875
+ $Y=0.0360 $X2=0.4070 $Y2=0.0360
r7 20 21 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3605
+ $Y=0.0360 $X2=0.3875 $Y2=0.0360
r8 19 20 7.92845 $w=1.3e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3265
+ $Y=0.0360 $X2=0.3605 $Y2=0.0360
r9 10 12 1.03257 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3085 $Y=0.0360 $X2=0.2970 $Y2=0.0360
r10 10 19 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3085
+ $Y=0.0360 $X2=0.3265 $Y2=0.0360
r11 12 18 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.2970 $Y2=0.0540
r12 9 17 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0720 $X2=0.2970 $Y2=0.0900
r13 9 18 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0720 $X2=0.2970 $Y2=0.0540
r14 16 17 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2835 $Y=0.0900 $X2=0.2970 $Y2=0.0900
r15 11 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0900 $X2=0.2835 $Y2=0.0900
r16 11 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0900
+ $X2=0.2700 $Y2=0.0945
r17 1 15 23.8708 $w=2.02e-08 $l=4.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.2700 $Y=0.0540 $X2=0.2700 $Y2=0.0945
r18 14 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r19 7 13 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r20 1 7 1e-05
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%PD1 VSS 12 13 29 8 2 9 7 1
c1 1 VSS 0.0035212f
c2 2 VSS 0.00387631f
c3 7 VSS 0.00288873f
c4 8 VSS 0.00232389f
c5 9 VSS 0.00245622f
r1 29 28 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.0675 $X2=0.6085 $Y2=0.0675
r2 27 28 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6040 $Y=0.0675 $X2=0.6085 $Y2=0.0675
r3 8 27 0.123457 $w=8.1e-08 $l=1e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.0675 $X2=0.6040 $Y2=0.0675
r4 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0675
+ $X2=0.5900 $Y2=0.0720
r5 23 24 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.5805
+ $Y=0.0720 $X2=0.5900 $Y2=0.0720
r6 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0720 $X2=0.5805 $Y2=0.0720
r7 21 22 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.0720 $X2=0.5670 $Y2=0.0720
r8 20 21 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0720 $X2=0.5400 $Y2=0.0720
r9 19 20 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5020
+ $Y=0.0720 $X2=0.5130 $Y2=0.0720
r10 18 19 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4805
+ $Y=0.0720 $X2=0.5020 $Y2=0.0720
r11 17 18 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.4540
+ $Y=0.0720 $X2=0.4805 $Y2=0.0720
r12 16 17 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4440
+ $Y=0.0720 $X2=0.4540 $Y2=0.0720
r13 15 16 1.63233 $w=1.3e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.4370
+ $Y=0.0720 $X2=0.4440 $Y2=0.0720
r14 14 15 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4280
+ $Y=0.0720 $X2=0.4370 $Y2=0.0720
r15 9 14 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4205
+ $Y=0.0720 $X2=0.4280 $Y2=0.0720
r16 1 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4280 $Y2=0.0720
r17 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r18 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r19 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0675 $X2=0.4320 $Y2=0.0675
r20 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4175 $Y2=0.0675
r21 2 8 1e-05
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%MH VSS 9 56 60 63 67 10 3 21 17 4 1 12 14 18 20
+ 16 19 15
c1 1 VSS 0.000220714f
c2 3 VSS 0.004653f
c3 4 VSS 0.00525505f
c4 9 VSS 0.0361288f
c5 10 VSS 0.00227891f
c6 11 VSS 0.000101038f
c7 12 VSS 0.00210173f
c8 13 VSS 6.81208e-20
c9 14 VSS 0.00869856f
c10 15 VSS 0.00780288f
c11 16 VSS 0.00150592f
c12 17 VSS 0.000570268f
c13 18 VSS 0.00101283f
c14 19 VSS 0.00309883f
c15 20 VSS 6.00843e-20
c16 21 VSS 0.00249794f
r1 67 66 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.2295 $X2=0.6085 $Y2=0.2295
r2 65 66 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6040 $Y=0.2295 $X2=0.6085 $Y2=0.2295
r3 3 65 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5920 $Y=0.2295 $X2=0.6040 $Y2=0.2295
r4 13 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2295 $X2=0.5920 $Y2=0.2295
r5 61 62 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.1890 $X2=0.5840 $Y2=0.1890
r6 63 61 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.1890 $X2=0.5795 $Y2=0.1890
r7 12 62 0.185185 $w=5.4e-08 $l=1e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.1890 $X2=0.5840 $Y2=0.1890
r8 12 3 0.518519 $w=3.9e-08 $l=4.05494e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.1890 $X2=0.5920 $Y2=0.2295
r9 60 59 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r10 58 59 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6580 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r11 4 58 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6460 $Y=0.0405 $X2=0.6580 $Y2=0.0405
r12 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0405 $X2=0.6460 $Y2=0.0405
r13 10 4 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0810 $X2=0.6460 $Y2=0.0810
r14 56 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.0810 $X2=0.6335 $Y2=0.0810
r15 3 48 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2295
+ $X2=0.5900 $Y2=0.2340
r16 4 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.0405
+ $X2=0.6440 $Y2=0.0360
r17 45 46 1.63233 $w=1.3e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.5990
+ $Y=0.2340 $X2=0.6060 $Y2=0.2340
r18 45 48 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5990
+ $Y=0.2340 $X2=0.5900 $Y2=0.2340
r19 44 46 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.6105
+ $Y=0.2340 $X2=0.6060 $Y2=0.2340
r20 43 44 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6305
+ $Y=0.2340 $X2=0.6105 $Y2=0.2340
r21 14 21 4.53042 $w=1.46981e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6665 $Y=0.2340 $X2=0.6930 $Y2=0.2340
r22 14 43 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.6665
+ $Y=0.2340 $X2=0.6305 $Y2=0.2340
r23 15 40 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.6530
+ $Y=0.0360 $X2=0.6705 $Y2=0.0360
r24 15 42 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6530
+ $Y=0.0360 $X2=0.6440 $Y2=0.0360
r25 21 39 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.2340 $X2=0.6930 $Y2=0.2160
r26 19 34 2.43171 $w=1.804e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6930 $Y=0.0360 $X2=0.6930 $Y2=0.0535
r27 19 40 3.59766 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.0360 $X2=0.6705 $Y2=0.0360
r28 38 39 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1980 $X2=0.6930 $Y2=0.2160
r29 37 38 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1800 $X2=0.6930 $Y2=0.1980
r30 36 37 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1680 $X2=0.6930 $Y2=0.1800
r31 35 36 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1590 $X2=0.6930 $Y2=0.1680
r32 17 20 2.43413 $w=1.59032e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6930 $Y=0.1465 $X2=0.6930 $Y2=0.1310
r33 17 35 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1465 $X2=0.6930 $Y2=0.1590
r34 33 34 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.0625 $X2=0.6930 $Y2=0.0535
r35 32 33 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.0720 $X2=0.6930 $Y2=0.0625
r36 31 32 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.0900 $X2=0.6930 $Y2=0.0720
r37 30 31 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1025 $X2=0.6930 $Y2=0.0900
r38 16 20 2.78392 $w=1.56471e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6930 $Y=0.1140 $X2=0.6930 $Y2=0.1310
r39 16 30 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1140 $X2=0.6930 $Y2=0.1025
r40 20 28 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1310 $X2=0.7110 $Y2=0.1310
r41 27 28 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1310 $X2=0.7110 $Y2=0.1310
r42 18 26 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.1310 $X2=0.7830 $Y2=0.1310
r43 18 27 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.1310 $X2=0.7290 $Y2=0.1310
r44 1 23 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.7830
+ $Y=0.1310 $X2=0.7830 $Y2=0.1310
r45 1 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7830 $Y=0.1310
+ $X2=0.7830 $Y2=0.1310
r46 9 23 0.314665 $w=2.27e-07 $l=4e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.7830 $Y=0.1350 $X2=0.7830 $Y2=0.1310
r47 3 12 1e-05
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%noxref_32 VSS 1
c1 1 VSS 0.00369864f
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%noxref_31 VSS 1
c1 1 VSS 0.00351511f
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%noxref_35 VSS 1
c1 1 VSS 0.00485788f
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%PD5 VSS 7 12 1 4 5
c1 1 VSS 0.00745215f
c2 4 VSS 0.00187448f
c3 5 VSS 0.00237127f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9890 $Y=0.0405 $X2=0.9865 $Y2=0.0405
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9740 $Y=0.0405 $X2=0.9865 $Y2=0.0405
r3 9 5 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.9585
+ $Y=0.0405 $X2=0.9720 $Y2=0.0405
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.9435
+ $Y=0.0405 $X2=0.9585 $Y2=0.0405
r5 1 8 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.9180
+ $Y=0.0405 $X2=0.9435 $Y2=0.0405
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9035 $Y=0.0405 $X2=0.9160 $Y2=0.0405
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9010 $Y=0.0405 $X2=0.9035 $Y2=0.0405
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%QN VSS 19 13 25 10 7 11 2 1 8 9
c1 1 VSS 0.00818693f
c2 2 VSS 0.00837846f
c3 7 VSS 0.00360063f
c4 8 VSS 0.0035953f
c5 9 VSS 0.00303755f
c6 10 VSS 0.00602154f
c7 11 VSS 0.00601229f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.2815 $Y=0.2025 $X2=1.2940 $Y2=0.2025
r2 25 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.2790 $Y=0.2025 $X2=1.2815 $Y2=0.2025
r3 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.2960 $Y=0.2025
+ $X2=1.2960 $Y2=0.2340
r4 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.2960
+ $Y=0.2340 $X2=1.3095 $Y2=0.2340
r5 11 20 1.09329 $w=1.76154e-08 $l=9.8e-09 $layer=M1 $thickness=3.6e-08
+ $X=1.3230 $Y=0.2340 $X2=1.3230 $Y2=0.2242
r6 11 23 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3230 $Y=0.2340 $X2=1.3095 $Y2=0.2340
r7 19 20 0.291487 $w=1.3e-08 $l=1.2e-09 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.2230 $X2=1.3230 $Y2=0.2242
r8 19 18 2.73998 $w=1.3e-08 $l=1.18e-08 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.2230 $X2=1.3230 $Y2=0.2112
r9 17 18 15.4488 $w=1.3e-08 $l=6.62e-08 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.1450 $X2=1.3230 $Y2=0.2112
r10 9 16 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3230 $Y=0.0675 $X2=1.3230 $Y2=0.0360
r11 9 17 18.0722 $w=1.3e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.0675 $X2=1.3230 $Y2=0.1450
r12 15 16 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3095 $Y=0.0360 $X2=1.3230 $Y2=0.0360
r13 14 15 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.2960
+ $Y=0.0360 $X2=1.3095 $Y2=0.0360
r14 10 14 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.2845
+ $Y=0.0360 $X2=1.2960 $Y2=0.0360
r15 1 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.2960 $Y=0.0675
+ $X2=1.2960 $Y2=0.0360
r16 7 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.2815 $Y=0.0675 $X2=1.2940 $Y2=0.0675
r17 13 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.2790 $Y=0.0675 $X2=1.2815 $Y2=0.0675
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%noxref_36 VSS 1
c1 1 VSS 0.00457305f
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%SEN VSS 9 45 50 3 4 13 14 1 15 11 12 10 16
c1 1 VSS 0.00392184f
c2 3 VSS 0.00899584f
c3 4 VSS 0.00830424f
c4 9 VSS 0.0816258f
c5 10 VSS 0.00452545f
c6 11 VSS 0.00483663f
c7 12 VSS 0.0016674f
c8 13 VSS 0.00325758f
c9 14 VSS 0.0008075f
c10 15 VSS 0.00610301f
c11 16 VSS 0.0117309f
r1 50 49 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.2050 $Y=0.2025 $X2=1.2025 $Y2=0.2025
r2 11 49 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.1900 $Y=0.2025 $X2=1.2025 $Y2=0.2025
r3 4 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.1880 $Y=0.2295
+ $X2=1.1880 $Y2=0.2340
r4 45 44 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.2050 $Y=0.0675 $X2=1.2025 $Y2=0.0675
r5 10 44 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.1900 $Y=0.0675 $X2=1.2025 $Y2=0.0675
r6 41 42 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.1745
+ $Y=0.2340 $X2=1.1880 $Y2=0.2340
r7 15 37 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1610 $Y=0.2340 $X2=1.1610 $Y2=0.2125
r8 15 41 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1610 $Y=0.2340 $X2=1.1745 $Y2=0.2340
r9 3 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.1725 $Y=0.0405
+ $X2=1.1610 $Y2=0.0515
r10 3 10 4.30736 $w=5.12e-08 $l=2.95e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.1725 $Y=0.0405 $X2=1.1725 $Y2=0.0700
r11 36 37 15.7403 $w=1.3e-08 $l=6.75e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.1450 $X2=1.1610 $Y2=0.2125
r12 35 36 14.9241 $w=1.3e-08 $l=6.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0810 $X2=1.1610 $Y2=0.1450
r13 34 35 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0650 $X2=1.1610 $Y2=0.0810
r14 33 34 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0515 $X2=1.1610 $Y2=0.0650
r15 32 33 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0425 $X2=1.1610 $Y2=0.0515
r16 13 32 1.28254 $w=1.3e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0370 $X2=1.1610 $Y2=0.0425
r17 30 35 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=1.1610 $Y=0.0810
+ $X2=1.1610 $Y2=0.0810
r18 29 30 27.2832 $w=1.3e-08 $l=1.17e-07 $layer=M2 $thickness=3.6e-08 $X=1.0440
+ $Y=0.0810 $X2=1.1610 $Y2=0.0810
r19 28 29 29.3819 $w=1.3e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.9180
+ $Y=0.0810 $X2=1.0440 $Y2=0.0810
r20 27 28 67.1587 $w=1.3e-08 $l=2.88e-07 $layer=M2 $thickness=3.6e-08 $X=0.6300
+ $Y=0.0810 $X2=0.9180 $Y2=0.0810
r21 26 27 65.0599 $w=1.3e-08 $l=2.79e-07 $layer=M2 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0810 $X2=0.6300 $Y2=0.0810
r22 16 26 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.3395
+ $Y=0.0810 $X2=0.3510 $Y2=0.0810
r23 14 22 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.0720 $X2=0.3510 $Y2=0.0855
r24 14 26 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.3510 $Y=0.0720 $X2=0.3510
+ $Y2=0.0810
r25 22 23 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0855 $X2=0.3510 $Y2=0.0945
r26 22 26 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.3510 $Y=0.0855 $X2=0.3510
+ $Y2=0.0810
r27 21 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1080 $X2=0.3510 $Y2=0.0945
r28 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1215 $X2=0.3510 $Y2=0.1080
r29 12 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1215
r30 9 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r31 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
r32 4 11 1e-05
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%SS VSS 9 34 39 13 15 14 17 16 12 3 4 1 11 10
c1 1 VSS 0.00110505f
c2 3 VSS 0.00589326f
c3 4 VSS 0.00659765f
c4 9 VSS 0.0384123f
c5 10 VSS 0.00326373f
c6 11 VSS 0.00339044f
c7 12 VSS 0.000970332f
c8 13 VSS 0.00841813f
c9 14 VSS 0.00177833f
c10 15 VSS 0.00265494f
c11 16 VSS 0.00614247f
c12 17 VSS 0.00201201f
r1 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0655 $Y=0.2295 $X2=1.0780 $Y2=0.2295
r2 39 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0630 $Y=0.2295 $X2=1.0655 $Y2=0.2295
r3 4 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0800 $Y=0.2295
+ $X2=1.0800 $Y2=0.2340
r4 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.0800
+ $Y=0.2340 $X2=1.0935 $Y2=0.2340
r5 16 32 7.21452 $w=1.425e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.2340 $X2=1.1070 $Y2=0.1980
r6 16 37 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1070 $Y=0.2340 $X2=1.0935 $Y2=0.2340
r7 10 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.0655 $Y=0.0405 $X2=1.0780 $Y2=0.0405
r8 34 10 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.0630 $Y=0.0405 $X2=1.0655 $Y2=0.0405
r9 31 32 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.1440 $X2=1.1070 $Y2=0.1980
r10 14 30 8.95608 $w=1.36627e-08 $l=4.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1070 $Y=0.0810 $X2=1.1070 $Y2=0.0395
r11 14 31 14.691 $w=1.3e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.0810 $X2=1.1070 $Y2=0.1440
r12 3 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0800 $Y=0.0405
+ $X2=1.0800 $Y2=0.0360
r13 17 29 1.40651 $w=1.51875e-08 $l=1.45774e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1070 $Y=0.0305 $X2=1.0935 $Y2=0.0360
r14 17 30 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.0305 $X2=1.1070 $Y2=0.0395
r15 28 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.0800
+ $Y=0.0360 $X2=1.0935 $Y2=0.0360
r16 27 28 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.0685
+ $Y=0.0360 $X2=1.0800 $Y2=0.0360
r17 26 27 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.0640
+ $Y=0.0360 $X2=1.0685 $Y2=0.0360
r18 25 26 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.0360 $X2=1.0640 $Y2=0.0360
r19 13 15 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0260 $Y=0.0360 $X2=0.9990 $Y2=0.0360
r20 13 25 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.0360 $X2=1.0530 $Y2=0.0360
r21 12 22 8.04505 $w=1.3e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.9990
+ $Y=0.0705 $X2=0.9990 $Y2=0.1050
r22 12 15 6.39593 $w=1.55565e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9990 $Y=0.0705 $X2=0.9990 $Y2=0.0360
r23 1 19 2.36633 $w=2.3e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.9990
+ $Y=0.1055 $X2=0.9990 $Y2=0.1055
r24 1 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.9990 $Y=0.1055
+ $X2=0.9990 $Y2=0.1050
r25 9 19 0.314665 $w=2.27e-07 $l=2.95e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.9990 $Y=0.1350 $X2=0.9990 $Y2=0.1055
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%MS VSS 10 43 46 51 53 3 15 12 13 1 17 4 11 18 19
+ 14 16
c1 1 VSS 0.00301528f
c2 3 VSS 0.00565664f
c3 4 VSS 0.00929567f
c4 10 VSS 0.0377166f
c5 11 VSS 0.00310098f
c6 12 VSS 0.00293078f
c7 13 VSS 0.00245475f
c8 14 VSS 0.00092433f
c9 15 VSS 0.00441658f
c10 16 VSS 0.00193943f
c11 17 VSS 0.000917797f
c12 18 VSS 0.00136404f
c13 19 VSS 0.00117518f
c14 20 VSS 0.00290094f
r1 53 52 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8810 $Y=0.2295 $X2=0.8785 $Y2=0.2295
r2 13 52 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8660 $Y=0.2295 $X2=0.8785 $Y2=0.2295
r3 12 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.2295 $X2=0.8080 $Y2=0.2295
r4 51 12 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.2295 $X2=0.7955 $Y2=0.2295
r5 48 13 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8370 $Y=0.2295 $X2=0.8640 $Y2=0.2295
r6 4 48 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08 $X=0.8100
+ $Y=0.2295 $X2=0.8370 $Y2=0.2295
r7 4 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8100 $Y=0.2295
+ $X2=0.8125 $Y2=0.2340
r8 15 20 4.06404 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8125 $Y=0.2340 $X2=0.8370 $Y2=0.2340
r9 46 45 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8270 $Y=0.0405 $X2=0.8245 $Y2=0.0405
r10 44 45 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8200 $Y=0.0405 $X2=0.8245 $Y2=0.0405
r11 3 44 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8080 $Y=0.0405 $X2=0.8200 $Y2=0.0405
r12 11 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.0405 $X2=0.8080 $Y2=0.0405
r13 43 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.0405 $X2=0.7955 $Y2=0.0405
r14 20 39 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.2340 $X2=0.8370 $Y2=0.2160
r15 3 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8100 $Y=0.0405
+ $X2=0.8100 $Y2=0.0535
r16 38 39 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1870 $X2=0.8370 $Y2=0.2160
r17 37 38 4.89699 $w=1.3e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1660 $X2=0.8370 $Y2=0.1870
r18 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1525 $X2=0.8370 $Y2=0.1660
r19 35 36 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1310 $X2=0.8370 $Y2=0.1525
r20 34 35 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1115 $X2=0.8370 $Y2=0.1310
r21 17 31 1.15159 $w=1.75e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1000 $X2=0.8370 $Y2=0.0900
r22 17 34 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1000 $X2=0.8370 $Y2=0.1115
r23 16 32 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0625 $X2=0.8100 $Y2=0.0720
r24 16 33 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0625 $X2=0.8100 $Y2=0.0535
r25 30 31 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8235 $Y=0.0900 $X2=0.8370 $Y2=0.0900
r26 19 28 1.38478 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.0900 $X2=0.7990 $Y2=0.0900
r27 19 30 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.0900 $X2=0.8235 $Y2=0.0900
r28 19 32 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0900 $X2=0.8100 $Y2=0.0720
r29 27 28 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.7765
+ $Y=0.0900 $X2=0.7990 $Y2=0.0900
r30 14 27 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.7470
+ $Y=0.0900 $X2=0.7765 $Y2=0.0900
r31 14 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7470 $Y=0.0900
+ $X2=0.7500 $Y2=0.0900
r32 14 18 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7470
+ $Y=0.0900 $X2=0.7290 $Y2=0.0900
r33 25 26 5.02115 $w=1.53e-08 $l=8.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.7415 $Y=0.0900 $X2=0.7500 $Y2=0.0900
r34 23 25 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.7385 $Y=0.0900 $X2=0.7415 $Y2=0.0900
r35 1 23 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.7285
+ $Y=0.0900 $X2=0.7385 $Y2=0.0900
r36 1 22 2.48102 $w=2.2e-08 $l=5e-10 $layer=LIG $thickness=4.8e-08 $X=0.7285
+ $Y=0.0900 $X2=0.7290 $Y2=0.0900
r37 22 25 1.47681 $w=1.53e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7290 $Y=0.0900 $X2=0.7415 $Y2=0.0900
r38 10 22 0.314665 $w=2.27e-07 $l=4.5e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.7290 $Y=0.1350 $X2=0.7290 $Y2=0.0900
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%SE VSS 34 5 6 9 13 8 12 1 2 10 7 11
c1 1 VSS 0.00197796f
c2 2 VSS 0.00380434f
c3 5 VSS 0.0426527f
c4 6 VSS 0.0802639f
c5 7 VSS 0.00172949f
c6 8 VSS 0.000586469f
c7 9 VSS 0.00475907f
c8 10 VSS 0.00582451f
c9 11 VSS 0.00128513f
c10 12 VSS 0.00721629f
c11 13 VSS 0.0561767f
r1 1 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
r2 5 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r3 38 39 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2745
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r4 37 38 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2595
+ $Y=0.1350 $X2=0.2745 $Y2=0.1350
r5 36 37 0.699569 $w=1.3e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.1350 $X2=0.2595 $Y2=0.1350
r6 34 8 2.49951 $w=7.46154e-09 $l=1.95256e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.1340 $X2=0.2445 $Y2=0.1350
r7 8 36 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2445
+ $Y=0.1350 $X2=0.2565 $Y2=0.1350
r8 34 11 0.433689 $w=1.8e-08 $l=4.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.1340 $X2=0.2250 $Y2=0.1297
r9 11 32 3.53073 $w=1.4087e-08 $l=1.72e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.1297 $X2=0.2250 $Y2=0.1125
r10 10 28 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.2250 $Y=0.0360 $X2=0.2250
+ $Y2=0.0450
r11 31 32 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0900 $X2=0.2250 $Y2=0.1125
r12 30 31 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0675 $X2=0.2250 $Y2=0.0900
r13 7 30 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0495 $X2=0.2250 $Y2=0.0675
r14 7 28 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.2250 $Y=0.0495 $X2=0.2250
+ $Y2=0.0450
r15 7 10 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.0495 $X2=0.2250 $Y2=0.0360
r16 28 29 14.108 $w=1.3e-08 $l=6.05e-08 $layer=M2 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0450 $X2=0.2855 $Y2=0.0450
r17 26 29 109.716 $w=1.3e-08 $l=4.705e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.7560 $Y=0.0450 $X2=0.2855 $Y2=0.0450
r18 13 24 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=1.1905
+ $Y=0.0450 $X2=1.2150 $Y2=0.0450
r19 13 26 101.321 $w=1.3e-08 $l=4.345e-07 $layer=M2 $thickness=3.6e-08
+ $X=1.1905 $Y=0.0450 $X2=0.7560 $Y2=0.0450
r20 12 24 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=1.2150 $Y=0.0360 $X2=1.2150
+ $Y2=0.0450
r21 20 21 6.41272 $w=1.3e-08 $l=2.75e-08 $layer=M1 $thickness=3.6e-08 $X=1.2150
+ $Y=0.1085 $X2=1.2150 $Y2=0.1360
r22 19 20 8.51143 $w=1.3e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=1.2150
+ $Y=0.0720 $X2=1.2150 $Y2=0.1085
r23 9 19 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.2150
+ $Y=0.0495 $X2=1.2150 $Y2=0.0720
r24 9 12 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.2150 $Y=0.0495 $X2=1.2150 $Y2=0.0360
r25 9 24 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=1.2150 $Y=0.0495 $X2=1.2150
+ $Y2=0.0450
r26 6 2 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=1.2150
+ $Y=0.1350 $X2=1.2150 $Y2=0.1360
r27 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.2150 $Y=0.1360
+ $X2=1.2150 $Y2=0.1360
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%SH VSS 11 12 65 68 70 73 14 25 21 23 6 13 18 16
+ 17 5 22 20 2 15 1 19 24
c1 1 VSS 0.00061553f
c2 2 VSS 0.0036769f
c3 5 VSS 0.0049921f
c4 6 VSS 0.00512208f
c5 11 VSS 0.037494f
c6 12 VSS 0.0801624f
c7 13 VSS 0.00374495f
c8 14 VSS 0.00392764f
c9 15 VSS 0.00818038f
c10 16 VSS 0.000578469f
c11 17 VSS 0.00138908f
c12 18 VSS 0.00125333f
c13 19 VSS 0.000144763f
c14 20 VSS 0.00335578f
c15 21 VSS 0.00649902f
c16 22 VSS 0.00215251f
c17 23 VSS 0.000116742f
c18 24 VSS 0.000366497f
c19 25 VSS 0.010681f
r1 73 72 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8810 $Y=0.0405 $X2=0.8785 $Y2=0.0405
r2 5 72 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8660 $Y=0.0405 $X2=0.8785 $Y2=0.0405
r3 69 5 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8540 $Y=0.0405 $X2=0.8660 $Y2=0.0405
r4 13 69 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.0405 $X2=0.8540 $Y2=0.0405
r5 70 13 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.0405 $X2=0.8495 $Y2=0.0405
r6 68 67 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9350 $Y=0.2295 $X2=0.9325 $Y2=0.2295
r7 66 67 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9280 $Y=0.2295 $X2=0.9325 $Y2=0.2295
r8 6 66 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9160 $Y=0.2295 $X2=0.9280 $Y2=0.2295
r9 14 6 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9035 $Y=0.2295 $X2=0.9160 $Y2=0.2295
r10 65 14 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9010 $Y=0.2295 $X2=0.9035 $Y2=0.2295
r11 5 57 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.0405
+ $X2=0.8640 $Y2=0.0360
r12 6 52 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.9180 $Y=0.2295
+ $X2=0.9180 $Y2=0.2340
r13 2 49 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.2690 $Y=0.1360
+ $X2=1.2690 $Y2=0.1445
r14 12 2 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=1.2690
+ $Y=0.1350 $X2=1.2690 $Y2=0.1360
r15 57 58 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.0360 $X2=0.8775 $Y2=0.0360
r16 55 58 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.0360 $X2=0.8775 $Y2=0.0360
r17 54 55 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.9020
+ $Y=0.0360 $X2=0.8910 $Y2=0.0360
r18 15 22 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.9200
+ $Y=0.0360 $X2=0.9450 $Y2=0.0360
r19 15 54 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.9200
+ $Y=0.0360 $X2=0.9020 $Y2=0.0360
r20 52 53 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.2340 $X2=0.9315 $Y2=0.2340
r21 21 53 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.2340 $X2=0.9315 $Y2=0.2340
r22 20 49 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.2690
+ $Y=0.1085 $X2=1.2690 $Y2=0.1445
r23 22 43 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.0360 $X2=0.9450 $Y2=0.0630
r24 17 38 6.50021 $w=1.33448e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.1980 $X2=0.9450 $Y2=0.1690
r25 17 21 7.21452 $w=1.425e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.1980 $X2=0.9450 $Y2=0.2340
r26 47 49 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=1.2690 $Y=0.1530
+ $X2=1.2690 $Y2=0.1445
r27 46 47 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=1.2445
+ $Y=0.1530 $X2=1.2690 $Y2=0.1530
r28 45 46 9.91056 $w=1.3e-08 $l=4.25e-08 $layer=M2 $thickness=3.6e-08 $X=1.2020
+ $Y=0.1530 $X2=1.2445 $Y2=0.1530
r29 44 45 32.0636 $w=1.3e-08 $l=1.375e-07 $layer=M2 $thickness=3.6e-08
+ $X=1.0645 $Y=0.1530 $X2=1.2020 $Y2=0.1530
r30 25 44 27.8662 $w=1.3e-08 $l=1.195e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.9450 $Y=0.1530 $X2=1.0645 $Y2=0.1530
r31 25 39 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.9450 $Y=0.1530 $X2=0.9450
+ $Y2=0.1485
r32 42 43 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.0900 $X2=0.9450 $Y2=0.0630
r33 41 42 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1000 $X2=0.9450 $Y2=0.0900
r34 40 41 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1100 $X2=0.9450 $Y2=0.1000
r35 16 39 3.96423 $w=1.3e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1315 $X2=0.9450 $Y2=0.1485
r36 16 40 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1315 $X2=0.9450 $Y2=0.1100
r37 37 38 0.4592 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1645 $X2=0.9450 $Y2=0.1690
r38 23 37 0.714311 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1575 $X2=0.9450 $Y2=0.1645
r39 23 39 1.50855 $w=1.55e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1575 $X2=0.9450 $Y2=0.1485
r40 23 25 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.9450 $Y=0.1575 $X2=0.9450
+ $Y2=0.1530
r41 36 38 4.4015 $w=1.35e-08 $l=2.78927e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9720 $Y=0.1620 $X2=0.9450 $Y2=0.1690
r42 35 36 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9990
+ $Y=0.1620 $X2=0.9720 $Y2=0.1620
r43 18 24 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0260 $Y=0.1620 $X2=1.0530 $Y2=0.1620
r44 18 35 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.1620 $X2=0.9990 $Y2=0.1620
r45 24 33 0.915974 $w=2.10182e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0530 $Y=0.1620 $X2=1.0530 $Y2=0.1510
r46 32 33 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1400 $X2=1.0530 $Y2=0.1510
r47 19 32 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1250 $X2=1.0530 $Y2=0.1400
r48 1 29 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=1.0530
+ $Y=0.1400 $X2=1.0530 $Y2=0.1400
r49 1 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.0530 $Y=0.1400
+ $X2=1.0530 $Y2=0.1400
r50 11 29 0.314665 $w=2.27e-07 $l=5e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.0530 $Y=0.1350 $X2=1.0530 $Y2=0.1400
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%CLKB VSS 11 12 61 63 13 22 16 5 19 15 6 20 14 17
+ 18 2 1 21
c1 1 VSS 0.000143777f
c2 2 VSS 0.000185014f
c3 5 VSS 0.00731696f
c4 6 VSS 0.00724595f
c5 11 VSS 0.00449088f
c6 12 VSS 0.00459975f
c7 13 VSS 0.00719777f
c8 14 VSS 0.00722479f
c9 15 VSS 0.00587187f
c10 16 VSS 0.00360098f
c11 17 VSS 0.000136224f
c12 18 VSS 0.000559923f
c13 19 VSS 0.00503928f
c14 20 VSS 0.00309804f
c15 21 VSS 0.000169373f
c16 22 VSS 0.0195593f
r1 14 6 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1600 $Y2=0.2160
r2 63 14 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r3 6 56 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r4 13 5 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1600 $Y2=0.0540
r5 61 13 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r6 56 57 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r7 15 56 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1505
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r8 5 53 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r9 20 49 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.1890 $Y2=0.2160
r10 20 57 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2340 $X2=0.1755 $Y2=0.2340
r11 53 54 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r12 19 44 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1890 $Y2=0.0630
r13 19 54 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1755 $Y2=0.0360
r14 1 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6210 $Y=0.1350
+ $X2=0.6210 $Y2=0.1395
r15 11 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1350
r16 48 49 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1980 $X2=0.1890 $Y2=0.2160
r17 47 48 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1765 $X2=0.1890 $Y2=0.1980
r18 46 47 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1630 $X2=0.1890 $Y2=0.1765
r19 45 46 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1530 $X2=0.1890 $Y2=0.1630
r20 43 44 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0900 $X2=0.1890 $Y2=0.0630
r21 42 43 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1100 $X2=0.1890 $Y2=0.0900
r22 16 42 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1325 $X2=0.1890 $Y2=0.1100
r23 16 45 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1325 $X2=0.1890 $Y2=0.1530
r24 21 39 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1620 $X2=0.6210 $Y2=0.1395
r25 21 33 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.6210 $Y=0.1620 $X2=0.6210
+ $Y2=0.1530
r26 17 39 5.47996 $w=1.3e-08 $l=2.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1160 $X2=0.6210 $Y2=0.1395
r27 37 38 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1530 $X2=0.2045 $Y2=0.1530
r28 37 45 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1890 $Y=0.1530
+ $X2=0.1890 $Y2=0.1530
r29 35 38 16.2067 $w=1.3e-08 $l=6.95e-08 $layer=M2 $thickness=3.6e-08 $X=0.2740
+ $Y=0.1530 $X2=0.2045 $Y2=0.1530
r30 33 34 15.2739 $w=1.3e-08 $l=6.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1530 $X2=0.6865 $Y2=0.1530
r31 33 39 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.6210 $Y=0.1530 $X2=0.6210
+ $Y2=0.1395
r32 32 33 34.1623 $w=1.3e-08 $l=1.465e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.4745 $Y=0.1530 $X2=0.6210 $Y2=0.1530
r33 32 35 46.7545 $w=1.3e-08 $l=2.005e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.4745 $Y=0.1530 $X2=0.2740 $Y2=0.1530
r34 22 31 18.3054 $w=1.3e-08 $l=7.85e-08 $layer=M2 $thickness=3.6e-08 $X=0.8125
+ $Y=0.1530 $X2=0.8910 $Y2=0.1530
r35 22 34 29.3819 $w=1.3e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.8125
+ $Y=0.1530 $X2=0.6865 $Y2=0.1530
r36 29 31 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.8910 $Y=0.1440
+ $X2=0.8910 $Y2=0.1530
r37 18 29 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1135 $X2=0.8910 $Y2=0.1440
r38 12 2 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.8910
+ $Y=0.1350 $X2=0.8910 $Y2=0.1350
r39 2 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8910 $Y=0.1350
+ $X2=0.8910 $Y2=0.1440
.ends

.subckt PM_SDFLx1_ASAP7_75t_R%CLKN VSS 16 17 18 19 20 101 103 30 27 26 31 8 33
+ 21 22 1 9 35 25 23 2 28 34 10 5 29 3 32 24
c1 1 VSS 0.00155782f
c2 2 VSS 0.000248279f
c3 3 VSS 5.59602e-20
c4 4 VSS 1e-36
c5 5 VSS 0.000279552f
c6 8 VSS 0.00776257f
c7 9 VSS 0.0080076f
c8 10 VSS 0.00384658f
c9 16 VSS 0.059277f
c10 17 VSS 0.00581222f
c11 18 VSS 0.00508682f
c12 19 VSS 0.00438505f
c13 20 VSS 0.00531307f
c14 21 VSS 0.00670317f
c15 22 VSS 0.00663444f
c16 23 VSS 0.00824526f
c17 24 VSS 0.00189728f
c18 25 VSS 0.00444664f
c19 26 VSS 0.00384712f
c20 27 VSS 0.00111484f
c21 28 VSS 0.00249598f
c22 29 VSS 0.00141031f
c23 30 VSS 0.0037822f
c24 31 VSS 0.00205933f
c25 32 VSS 0.00401181f
c26 33 VSS 0.00139689f
c27 34 VSS 0.000675209f
c28 35 VSS 0.0312055f
r1 103 102 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r2 22 102 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r3 101 100 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r4 21 100 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r5 9 98 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0550 $Y2=0.2340
r6 8 95 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0550 $Y2=0.0360
r7 97 98 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.2340 $X2=0.0550 $Y2=0.2340
r8 26 97 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0460 $Y2=0.2340
r9 26 32 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0180 $Y2=0.2340
r10 94 95 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.0360 $X2=0.0550 $Y2=0.0360
r11 25 94 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0460 $Y2=0.0360
r12 25 30 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0180 $Y2=0.0360
r13 32 92 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.2340 $X2=0.0180 $Y2=0.2160
r14 30 91 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.0360 $X2=0.0180 $Y2=0.0630
r15 1 83 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
r16 16 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r17 24 31 1.81469 $w=1.6125e-08 $l=1.35831e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.2025 $X2=0.0165 $Y2=0.1890
r18 24 92 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.2025 $X2=0.0180 $Y2=0.2160
r19 90 91 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0900 $X2=0.0180 $Y2=0.0630
r20 89 90 9.67737 $w=1.3e-08 $l=4.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1315 $X2=0.0180 $Y2=0.0900
r21 23 31 2.63085 $w=1.54194e-08 $l=1.7066e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1720 $X2=0.0165 $Y2=0.1890
r22 23 89 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1720 $X2=0.0180 $Y2=0.1315
r23 2 74 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1355
+ $X2=0.5670 $Y2=0.1350
r24 17 2 3.19489 $w=1.24e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1355
r25 33 69 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.1350 $Y=0.1980 $X2=0.1350
+ $Y2=0.1890
r26 83 84 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1540
r27 81 84 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1720 $X2=0.1350 $Y2=0.1540
r28 27 69 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.1350 $Y=0.1845 $X2=0.1350
+ $Y2=0.1890
r29 27 81 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1845 $X2=0.1350 $Y2=0.1720
r30 27 33 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1845 $X2=0.1350 $Y2=0.1980
r31 78 79 1.90199 $w=1.38333e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.0255 $Y=0.1890 $X2=0.0345 $Y2=0.1890
r32 31 78 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0165
+ $Y=0.1890 $X2=0.0255 $Y2=0.1890
r33 34 71 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.1980 $X2=0.5670 $Y2=0.1845
r34 34 62 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.5670 $Y=0.1980 $X2=0.5670
+ $Y2=0.1890
r35 74 75 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1485
r36 72 75 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1620 $X2=0.5670 $Y2=0.1485
r37 28 71 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1755 $X2=0.5670 $Y2=0.1845
r38 28 72 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1755 $X2=0.5670 $Y2=0.1620
r39 69 70 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1890 $X2=0.1595 $Y2=0.1890
r40 68 69 11.8927 $w=1.3e-08 $l=5.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.0840
+ $Y=0.1890 $X2=0.1350 $Y2=0.1890
r41 67 68 11.8927 $w=1.3e-08 $l=5.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.0330
+ $Y=0.1890 $X2=0.0840 $Y2=0.1890
r42 67 79 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.0330 $Y=0.1890
+ $X2=0.0345 $Y2=0.1890
r43 63 64 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.6480
+ $Y=0.1890 $X2=0.7290 $Y2=0.1890
r44 62 63 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1890 $X2=0.6480 $Y2=0.1890
r45 62 71 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.5670 $Y=0.1890 $X2=0.5670
+ $Y2=0.1845
r46 35 62 46.7546 $w=1.3e-08 $l=2.005e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.3665 $Y=0.1890 $X2=0.5670 $Y2=0.1890
r47 35 70 48.2703 $w=1.3e-08 $l=2.07e-07 $layer=M2 $thickness=3.6e-08 $X=0.3665
+ $Y=0.1890 $X2=0.1595 $Y2=0.1890
r48 5 59 2.78395 $w=2.4e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.9450
+ $Y=0.1780 $X2=0.9450 $Y2=0.1780
r49 20 5 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.9450 $Y=0.1350 $X2=0.9450 $Y2=0.1780
r50 3 52 2.78395 $w=2.4e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.6750
+ $Y=0.1780 $X2=0.6750 $Y2=0.1780
r51 18 3 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.6750 $Y=0.1350 $X2=0.6750 $Y2=0.1780
r52 60 64 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.7290 $Y=0.1845
+ $X2=0.7290 $Y2=0.1890
r53 29 60 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1680 $X2=0.7290 $Y2=0.1845
r54 58 59 6.83711 $w=2.22e-08 $l=1.5e-09 $layer=LISD $thickness=2.7e-08
+ $X=0.9435 $Y=0.1780 $X2=0.9450 $Y2=0.1780
r55 57 58 12.9145 $w=2.22e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9180 $Y=0.1780 $X2=0.9435 $Y2=0.1780
r56 56 57 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9045 $Y=0.1780 $X2=0.9180 $Y2=0.1780
r57 55 56 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8910 $Y=0.1780 $X2=0.9045 $Y2=0.1780
r58 54 55 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8775 $Y=0.1780 $X2=0.8910 $Y2=0.1780
r59 53 54 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8640 $Y=0.1780 $X2=0.8775 $Y2=0.1780
r60 51 52 12.9145 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6885 $Y=0.1780 $X2=0.6750 $Y2=0.1780
r61 50 51 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7155 $Y=0.1780 $X2=0.6885 $Y2=0.1780
r62 48 49 6.07743 $w=2.22e-08 $l=1.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7290 $Y=0.1780 $X2=0.7410 $Y2=0.1780
r63 48 60 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7290 $Y=0.1780
+ $X2=0.7290 $Y2=0.1845
r64 47 48 5.31775 $w=2.22e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7185 $Y=0.1780 $X2=0.7290 $Y2=0.1780
r65 47 50 1.51936 $w=2.22e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.7185
+ $Y=0.1780 $X2=0.7155 $Y2=0.1780
r66 46 49 4.55807 $w=2.22e-08 $l=9e-09 $layer=LISD $thickness=2.7e-08 $X=0.7500
+ $Y=0.1780 $X2=0.7410 $Y2=0.1780
r67 45 46 6.07743 $w=2.22e-08 $l=1.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7620 $Y=0.1780 $X2=0.7500 $Y2=0.1780
r68 44 45 4.05162 $w=2.22e-08 $l=8e-09 $layer=LISD $thickness=2.7e-08 $X=0.7700
+ $Y=0.1780 $X2=0.7620 $Y2=0.1780
r69 43 44 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7835 $Y=0.1780 $X2=0.7700 $Y2=0.1780
r70 42 43 6.58388 $w=2.22e-08 $l=1.3e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7965 $Y=0.1780 $X2=0.7835 $Y2=0.1780
r71 41 42 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8100 $Y=0.1780 $X2=0.7965 $Y2=0.1780
r72 10 41 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8370 $Y=0.1780 $X2=0.8100 $Y2=0.1780
r73 10 53 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8370 $Y=0.1780 $X2=0.8640 $Y2=0.1780
r74 4 40 2.78395 $w=2.4e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.8370
+ $Y=0.1780 $X2=0.8370 $Y2=0.1780
r75 4 10 10.3807 $w=2.30357e-08 $l=0 $layer=LISD $thickness=3.675e-08 $X=0.8370
+ $Y=0.1780 $X2=0.8370 $Y2=0.1780
r76 19 40 0.314665 $w=2.27e-07 $l=4.3e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.8370 $Y=0.1350 $X2=0.8370 $Y2=0.1780
r77 9 22 1e-05
r78 8 21 1e-05
.ends


*
.SUBCKT SDFLx1_ASAP7_75t_R VSS VDD CLK SE D SI QN
*
* VSS VSS
* VDD VDD
* CLK CLK
* SE SE
* D D
* SI SI
* QN QN
*
*

MM20 N_MM20_d N_MM20_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM23 N_MM23_d N_MM22_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM26 N_MM26_d N_MM31_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM29 N_MM29_d N_MM27_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM32 N_MM32_d N_MM30_g N_MM32_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM3_g N_MM5_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM10_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM6 N_MM6_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM12 N_MM12_d N_MM12_g N_MM12_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM17 N_MM17_d N_MM17_g N_MM17_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM16 N_MM16_d N_MM16_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM14 N_MM14_d N_MM14_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM0 N_MM0_d N_MM0_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24 N_MM24_d N_MM24_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM21 N_MM21_d N_MM20_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM22 N_MM22_d N_MM22_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM31 N_MM31_d N_MM31_g N_MM31_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM27 N_MM27_d N_MM27_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM30 N_MM30_d N_MM30_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g N_MM3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM13 N_MM13_d N_MM17_g N_MM13_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM18 N_MM18_d N_MM18_g N_MM18_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM19 N_MM19_d N_MM16_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM15 N_MM15_d N_MM14_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM2 N_MM2_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25 N_MM25_d N_MM24_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "SDFLx1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "SDFLx1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_SDFLx1_ASAP7_75t_R%NET0167 VSS N_MM29_d N_MM32_s N_NET0167_1
+ PM_SDFLx1_ASAP7_75t_R%NET0167
cc_1 N_NET0167_1 N_MM27_g 0.0172747f
cc_2 N_NET0167_1 N_MM30_g 0.0173178f
x_PM_SDFLx1_ASAP7_75t_R%NET0144 VSS N_MM31_s N_MM27_d N_MM30_d N_MM3_s
+ N_NET0144_9 N_NET0144_7 N_NET0144_1 N_NET0144_8 N_NET0144_2
+ PM_SDFLx1_ASAP7_75t_R%NET0144
cc_3 N_NET0144_9 N_CLKN_35 0.00293384f
cc_4 N_NET0144_7 N_SE_1 0.00103669f
cc_5 N_NET0144_9 N_SE_8 0.000722908f
cc_6 N_NET0144_1 N_MM31_g 0.000818607f
cc_7 N_NET0144_7 N_MM31_g 0.0328701f
cc_8 N_NET0144_7 N_SEN_1 0.000888104f
cc_9 N_NET0144_1 N_MM27_g 0.000832514f
cc_10 N_NET0144_9 N_SEN_12 0.00206291f
cc_11 N_NET0144_7 N_MM27_g 0.0329847f
cc_12 N_NET0144_8 N_D_1 0.000763936f
cc_13 N_NET0144_2 N_MM30_g 0.000895522f
cc_14 N_NET0144_9 N_D 0.00223149f
cc_15 N_NET0144_8 N_MM30_g 0.0332853f
cc_16 N_NET0144_9 N_SI_4 0.000664488f
cc_17 N_NET0144_2 N_MM3_g 0.000855506f
cc_18 N_NET0144_8 N_SI_1 0.000864798f
cc_19 N_NET0144_8 N_MM3_g 0.0335016f
cc_20 N_NET0144_7 N_PU1_11 0.000549395f
cc_21 N_NET0144_8 N_PU1_9 0.00110376f
cc_22 N_NET0144_7 N_PU1_8 0.000553928f
cc_23 N_NET0144_1 N_PU1_11 0.000608137f
cc_24 N_NET0144_8 N_PU1_2 0.00130938f
cc_25 N_NET0144_2 N_PU1_2 0.00160191f
cc_26 N_NET0144_1 N_PU1_1 0.00303674f
cc_27 N_NET0144_9 N_PU1_11 0.0126831f
x_PM_SDFLx1_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_SDFLx1_ASAP7_75t_R%noxref_24
cc_28 N_noxref_24_1 N_MM20_g 0.00368873f
cc_29 N_noxref_24_1 N_CLKN_31 3.33509e-20
cc_30 N_noxref_24_1 N_CLKN_8 0.000550469f
cc_31 N_noxref_24_1 N_CLKN_9 4.50378e-20
cc_32 N_noxref_24_1 N_CLKN_30 5.73411e-20
cc_33 N_noxref_24_1 N_CLKN_23 0.000387378f
cc_34 N_noxref_24_1 N_CLKN_21 0.0275999f
x_PM_SDFLx1_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_SDFLx1_ASAP7_75t_R%noxref_25
cc_35 N_noxref_25_1 N_MM20_g 0.00368306f
cc_36 N_noxref_25_1 N_CLKN_9 0.000467847f
cc_37 N_noxref_25_1 N_CLKN_8 4.3136e-20
cc_38 N_noxref_25_1 N_CLKN_32 5.34043e-20
cc_39 N_noxref_25_1 N_CLKN_24 7.85693e-20
cc_40 N_noxref_25_1 N_CLKN_31 9.41135e-20
cc_41 N_noxref_25_1 N_CLKN_23 0.000274533f
cc_42 N_noxref_25_1 N_CLKN_22 0.027668f
cc_43 N_noxref_25_1 N_noxref_24_1 0.00204688f
x_PM_SDFLx1_ASAP7_75t_R%noxref_30 VSS N_noxref_30_1
+ PM_SDFLx1_ASAP7_75t_R%noxref_30
cc_44 N_noxref_30_1 N_CLKN_2 0.000194373f
cc_45 N_noxref_30_1 N_MM1_g 0.0107895f
cc_46 N_noxref_30_1 N_MM3_g 0.00149853f
cc_47 N_noxref_30_1 N_SI_1 0.00278437f
cc_48 N_noxref_30_1 N_PU1_2 0.00114378f
cc_49 N_noxref_30_1 N_PU1_9 0.0161574f
cc_50 N_noxref_30_1 N_PU1_10 0.0551754f
cc_51 N_noxref_30_1 N_NET0168_8 0.0368029f
x_PM_SDFLx1_ASAP7_75t_R%PD4 VSS N_MM18_s N_MM19_d N_PD4_1
+ PM_SDFLx1_ASAP7_75t_R%PD4
cc_52 N_PD4_1 N_MM18_g 0.00776292f
cc_53 N_PD4_1 N_MM16_g 0.00781368f
x_PM_SDFLx1_ASAP7_75t_R%PD3 VSS N_MM9_s N_MM8_d N_PD3_1
+ PM_SDFLx1_ASAP7_75t_R%PD3
cc_54 N_PD3_1 N_MM9_g 0.00775919f
cc_55 N_PD3_1 N_MM11_g 0.00785068f
x_PM_SDFLx1_ASAP7_75t_R%PD2 VSS N_MM10_s N_MM11_d N_PD2_5 N_PD2_1 N_PD2_4
+ PM_SDFLx1_ASAP7_75t_R%PD2
cc_56 N_PD2_5 N_CLKN_29 8.73123e-20
cc_57 N_PD2_5 N_CLKN_10 0.0018237f
cc_58 N_PD2_5 N_CLKN_3 0.000276686f
cc_59 N_PD2_1 N_MM9_g 0.00205987f
cc_60 N_PD2_4 N_MM9_g 0.00712351f
cc_61 N_PD2_5 N_MM9_g 0.0239108f
cc_62 N_PD2_4 N_MM10_g 0.0150985f
cc_63 N_PD2_5 N_MM11_g 0.0146992f
cc_64 N_PD2_4 N_MH_14 0.000323301f
cc_65 N_PD2_1 N_MH_17 0.000362771f
cc_66 N_PD2_4 N_MH_3 0.000613285f
cc_67 N_PD2_1 N_MH_14 0.00311186f
x_PM_SDFLx1_ASAP7_75t_R%CLK VSS CLK N_MM20_g N_CLK_4 N_CLK_6 N_CLK_1 N_CLK_5
+ PM_SDFLx1_ASAP7_75t_R%CLK
x_PM_SDFLx1_ASAP7_75t_R%noxref_34 VSS N_noxref_34_1
+ PM_SDFLx1_ASAP7_75t_R%noxref_34
cc_68 N_noxref_34_1 N_MM0_g 0.00135211f
cc_69 N_noxref_34_1 N_SEN_3 0.000119668f
cc_70 N_noxref_34_1 N_SEN_4 0.000412374f
cc_71 N_noxref_34_1 N_SEN_11 0.0373001f
cc_72 N_noxref_34_1 N_noxref_31_1 0.000462467f
cc_73 N_noxref_34_1 N_noxref_32_1 0.00774935f
cc_74 N_noxref_34_1 N_noxref_33_1 0.00120774f
x_PM_SDFLx1_ASAP7_75t_R%noxref_33 VSS N_noxref_33_1
+ PM_SDFLx1_ASAP7_75t_R%noxref_33
cc_75 N_noxref_33_1 N_MM0_g 0.0013111f
cc_76 N_noxref_33_1 N_SEN_3 0.00191288f
cc_77 N_noxref_33_1 N_SEN_10 0.0378042f
cc_78 N_noxref_33_1 N_noxref_31_1 0.00744269f
cc_79 N_noxref_33_1 N_noxref_32_1 0.000450527f
x_PM_SDFLx1_ASAP7_75t_R%PU1 VSS N_MM31_d N_MM3_d N_MM1_s N_PU1_10 N_PU1_2
+ N_PU1_11 N_PU1_8 N_PU1_1 N_PU1_9 PM_SDFLx1_ASAP7_75t_R%PU1
cc_80 N_PU1_10 N_CLKN_28 0.000377961f
cc_81 N_PU1_10 N_MM22_g 3.23234e-20
cc_82 N_PU1_10 N_CLKN_35 8.12706e-20
cc_83 N_PU1_10 N_CLKN_2 0.00104401f
cc_84 N_PU1_10 N_CLKN_34 0.000367896f
cc_85 N_PU1_2 N_MM1_g 0.0015956f
cc_86 N_PU1_11 N_CLKN_35 0.00328784f
cc_87 N_PU1_10 N_MM1_g 0.033968f
cc_88 N_PU1_8 N_SE_8 0.000736071f
cc_89 N_PU1_8 N_SE_1 0.00101689f
cc_90 N_PU1_1 N_MM31_g 0.00131787f
cc_91 N_PU1_8 N_MM31_g 0.0341707f
cc_92 N_PU1_2 N_SI_5 0.000617683f
cc_93 N_PU1_9 N_SI_1 0.00196303f
cc_94 N_PU1_2 N_SI_6 0.00293934f
cc_95 N_PU1_11 N_SI_6 0.00310512f
cc_96 N_PU1_9 N_MM3_g 0.0347119f
cc_97 N_PU1_2 N_MH_3 0.00118746f
cc_98 N_PU1_2 N_MH_12 0.00293214f
x_PM_SDFLx1_ASAP7_75t_R%noxref_27 VSS N_noxref_27_1
+ PM_SDFLx1_ASAP7_75t_R%noxref_27
cc_99 N_noxref_27_1 N_CLKN_1 0.000138589f
cc_100 N_noxref_27_1 N_MM22_g 0.00341439f
cc_101 N_noxref_27_1 N_CLKB_6 0.000367294f
cc_102 N_noxref_27_1 N_CLKB_14 0.0271182f
cc_103 N_noxref_27_1 N_PU1_8 0.000585889f
cc_104 N_noxref_27_1 N_noxref_26_1 0.00148647f
x_PM_SDFLx1_ASAP7_75t_R%noxref_29 VSS N_noxref_29_1
+ PM_SDFLx1_ASAP7_75t_R%noxref_29
cc_105 N_noxref_29_1 N_MM31_g 0.00147824f
cc_106 N_noxref_29_1 N_CLKB_14 0.000652468f
cc_107 N_noxref_29_1 N_PU1_8 0.0361347f
cc_108 N_noxref_29_1 N_noxref_26_1 0.00046969f
cc_109 N_noxref_29_1 N_noxref_27_1 0.00770807f
cc_110 N_noxref_29_1 N_noxref_28_1 0.00123606f
x_PM_SDFLx1_ASAP7_75t_R%noxref_28 VSS N_noxref_28_1
+ PM_SDFLx1_ASAP7_75t_R%noxref_28
cc_111 N_noxref_28_1 N_MM31_g 0.00163805f
cc_112 N_noxref_28_1 N_CLKB_13 0.000604377f
cc_113 N_noxref_28_1 N_NET0168_7 0.0361899f
cc_114 N_noxref_28_1 N_noxref_26_1 0.00770687f
cc_115 N_noxref_28_1 N_noxref_27_1 0.000469905f
x_PM_SDFLx1_ASAP7_75t_R%D VSS D N_MM30_g N_D_1 N_D_5 PM_SDFLx1_ASAP7_75t_R%D
cc_116 N_MM30_g N_SEN_16 0.000478536f
cc_117 N_MM30_g N_SEN_1 0.000814048f
cc_118 N_D_1 N_SEN_1 0.00132218f
cc_119 N_D_5 N_SEN_14 0.00179044f
cc_120 N_D N_SEN_12 0.00197214f
cc_121 N_MM30_g N_MM27_g 0.00504428f
x_PM_SDFLx1_ASAP7_75t_R%noxref_26 VSS N_noxref_26_1
+ PM_SDFLx1_ASAP7_75t_R%noxref_26
cc_122 N_noxref_26_1 N_CLKN_1 0.000144352f
cc_123 N_noxref_26_1 N_MM22_g 0.00338509f
cc_124 N_noxref_26_1 N_CLKB_5 0.000432383f
cc_125 N_noxref_26_1 N_CLKB_13 0.0270762f
cc_126 N_noxref_26_1 N_NET0168_7 0.000558204f
x_PM_SDFLx1_ASAP7_75t_R%SI VSS SI N_MM3_g N_SI_5 N_SI_6 N_SI_7 N_SI_4 N_SI_1
+ PM_SDFLx1_ASAP7_75t_R%SI
cc_127 N_SI_5 N_MM1_g 7.3915e-20
cc_128 N_SI_5 N_CLKN_2 0.00058192f
cc_129 N_SI_5 N_CLKN_35 0.00104747f
cc_130 N_SI_6 N_CLKN_35 0.000321682f
cc_131 N_SI_7 N_CLKN_28 0.000860886f
cc_132 N_SI_6 N_CLKN_34 0.000882831f
cc_133 N_SI_5 N_CLKN_28 0.00241179f
cc_134 N_SI_4 N_MM30_g 0.000933337f
cc_135 N_SI_1 N_D_1 0.000979599f
cc_136 N_MM3_g N_MM30_g 0.0040652f
x_PM_SDFLx1_ASAP7_75t_R%NET0168 VSS N_MM26_d N_MM5_s N_NET0168_7 N_NET0168_9
+ N_NET0168_1 N_NET0168_11 N_NET0168_12 N_NET0168_10 N_NET0168_2 N_NET0168_8
+ PM_SDFLx1_ASAP7_75t_R%NET0168
cc_137 N_NET0168_7 N_SE_1 0.00129827f
cc_138 N_NET0168_9 N_SE_10 0.000661871f
cc_139 N_NET0168_1 N_SE_8 0.000831645f
cc_140 N_NET0168_11 N_SE_7 0.00129296f
cc_141 N_NET0168_12 N_SE_10 0.00131306f
cc_142 N_NET0168_1 N_MM31_g 0.00154571f
cc_143 N_NET0168_11 N_SE_8 0.00362626f
cc_144 N_NET0168_10 N_SE_13 0.00427199f
cc_145 N_NET0168_7 N_MM31_g 0.034186f
cc_146 N_NET0168_10 N_SEN_12 0.000320068f
cc_147 N_NET0168_10 N_SEN_16 0.000390465f
cc_148 N_NET0168_11 N_SEN_12 0.00112606f
cc_149 N_NET0168_10 N_SEN_14 0.00530239f
cc_150 N_NET0168_2 N_MM3_g 0.00150903f
cc_151 N_NET0168_8 N_SI_1 0.00162109f
cc_152 N_NET0168_8 N_MM3_g 0.0345523f
x_PM_SDFLx1_ASAP7_75t_R%PD1 VSS N_MM32_d N_MM5_d N_MM4_s N_PD1_8 N_PD1_2
+ N_PD1_9 N_PD1_7 N_PD1_1 PM_SDFLx1_ASAP7_75t_R%PD1
cc_153 N_PD1_8 N_CLKN_28 0.000152897f
cc_154 N_PD1_8 N_CLKN_2 0.00113259f
cc_155 N_PD1_2 N_MM1_g 0.0011547f
cc_156 N_PD1_9 N_CLKN_28 0.00234083f
cc_157 N_PD1_8 N_MM1_g 0.0357125f
cc_158 N_PD1_9 N_SE_13 0.00220483f
cc_159 N_PD1_9 N_SEN_12 9.83162e-20
cc_160 N_PD1_9 N_MM27_g 0.000309102f
cc_161 N_PD1_9 N_SEN_14 0.000560625f
cc_162 N_PD1_9 N_SEN_16 0.00391671f
cc_163 N_PD1_7 N_D_1 0.000894761f
cc_164 N_PD1_1 N_MM30_g 0.00127495f
cc_165 N_PD1_9 N_D_5 0.00274403f
cc_166 N_PD1_7 N_MM30_g 0.0342193f
cc_167 N_PD1_1 N_MM3_g 0.000766737f
cc_168 N_PD1_7 N_SI_1 0.000891996f
cc_169 N_PD1_9 N_SI_7 0.00254764f
cc_170 N_PD1_7 N_MM3_g 0.0340534f
cc_171 N_PD1_8 N_CLKB_1 0.000985053f
cc_172 N_PD1_9 N_CLKB_17 0.00071161f
cc_173 N_PD1_2 N_MM10_g 0.000889176f
cc_174 N_PD1_9 N_CLKB_22 0.00090233f
cc_175 N_PD1_8 N_MM10_g 0.0329238f
cc_176 N_PD1_8 N_MH_10 0.00114164f
cc_177 N_PD1_9 N_MH_15 0.000953028f
cc_178 N_PD1_2 N_MH_4 0.00367285f
cc_179 N_PD1_7 N_NET0168_10 0.000584303f
cc_180 N_PD1_7 N_NET0168_8 0.00064714f
cc_181 N_PD1_9 N_NET0168_2 0.00066923f
cc_182 N_PD1_1 N_NET0168_2 0.00377826f
cc_183 N_PD1_9 N_NET0168_10 0.00913245f
x_PM_SDFLx1_ASAP7_75t_R%MH VSS N_MM7_g N_MM4_d N_MM9_d N_MM1_d N_MM10_d N_MH_10
+ N_MH_3 N_MH_21 N_MH_17 N_MH_4 N_MH_1 N_MH_12 N_MH_14 N_MH_18 N_MH_20 N_MH_16
+ N_MH_19 N_MH_15 PM_SDFLx1_ASAP7_75t_R%MH
cc_184 N_MH_10 N_CLKN_28 0.000126639f
cc_185 N_MH_10 N_CLKN_29 0.000348814f
cc_186 N_MH_10 N_MM1_g 0.000401025f
cc_187 N_MH_10 N_CLKN_2 0.000206389f
cc_188 N_MH_3 N_CLKN_34 0.000325817f
cc_189 N_MH_3 N_CLKN_28 0.000335674f
cc_190 N_MH_21 N_CLKN_29 0.000419151f
cc_191 N_MH_17 N_CLKN_29 0.00644609f
cc_192 N_MH_17 N_CLKN_3 0.000496837f
cc_193 N_MH_4 N_MM9_g 0.000618766f
cc_194 N_MH_1 N_CLKN_10 0.00215012f
cc_195 N_MH_12 N_CLKN_2 0.000666875f
cc_196 N_MH_17 N_CLKN_10 0.000744646f
cc_197 N_MH_14 N_CLKN_35 0.00140167f
cc_198 N_MH_18 N_CLKN_29 0.00150465f
cc_199 N_MH_3 N_MM1_g 0.00158418f
cc_200 N_MH_14 N_CLKN_34 0.00379103f
cc_201 N_MM7_g N_CLKN_10 0.00512105f
cc_202 N_MH_12 N_MM1_g 0.0329535f
cc_203 N_MM7_g N_MM12_g 0.0127127f
cc_204 N_MH_10 N_MM9_g 0.0361151f
cc_205 N_MH_10 N_CLKB_2 9.73291e-20
cc_206 N_MH_10 N_CLKB_17 0.000270079f
cc_207 N_MH_10 N_MM17_g 0.000141858f
cc_208 N_MH_3 N_CLKB_21 0.000304961f
cc_209 N_MH_20 N_CLKB_21 0.000316788f
cc_210 N_MH_14 N_CLKB_21 0.000452324f
cc_211 N_MH_12 N_MM10_g 0.0163577f
cc_212 N_MH_16 N_CLKB_17 0.000545553f
cc_213 N_MH_3 N_CLKB_1 0.000608409f
cc_214 N_MH_4 N_CLKB_17 0.0007682f
cc_215 N_MH_4 N_MM10_g 0.00113649f
cc_216 N_MH_3 N_MM10_g 0.00122003f
cc_217 N_MH_10 N_CLKB_1 0.00170375f
cc_218 N_MH_17 N_CLKB_21 0.00202765f
cc_219 N_MH_18 N_CLKB_22 0.0025362f
cc_220 N_MH_10 N_MM10_g 0.0527851f
cc_221 N_MH_19 N_MS_18 0.000280987f
cc_222 N_MH_4 N_MS_1 0.000395404f
cc_223 N_MH_18 N_MS_19 0.000419258f
cc_224 N_MH_18 N_MS_1 0.000673484f
cc_225 N_MM7_g N_MS_3 0.000958346f
cc_226 N_MH_1 N_MS_14 0.000962086f
cc_227 N_MH_18 N_MS_17 0.0010047f
cc_228 N_MH_1 N_MS_1 0.00130888f
cc_229 N_MM7_g N_MS_1 0.00223179f
cc_230 N_MM7_g N_MS_11 0.00638226f
cc_231 N_MM7_g N_MS_12 0.0064202f
cc_232 N_MH_16 N_MS_18 0.00432186f
cc_233 N_MH_18 N_MS_14 0.00561616f
cc_234 N_MM7_g N_MM11_g 0.0293989f
x_PM_SDFLx1_ASAP7_75t_R%noxref_32 VSS N_noxref_32_1
+ PM_SDFLx1_ASAP7_75t_R%noxref_32
cc_235 N_noxref_32_1 N_SEN_4 0.000149883f
cc_236 N_noxref_32_1 N_SEN_11 0.000881497f
cc_237 N_noxref_32_1 N_SS_11 0.01695f
cc_238 N_noxref_32_1 N_MM14_g 0.00579455f
cc_239 N_noxref_32_1 N_noxref_31_1 0.0015183f
x_PM_SDFLx1_ASAP7_75t_R%noxref_31 VSS N_noxref_31_1
+ PM_SDFLx1_ASAP7_75t_R%noxref_31
cc_240 N_noxref_31_1 N_SEN_3 0.00180026f
cc_241 N_noxref_31_1 N_SS_10 0.0168959f
cc_242 N_noxref_31_1 N_MM14_g 0.00570942f
x_PM_SDFLx1_ASAP7_75t_R%noxref_35 VSS N_noxref_35_1
+ PM_SDFLx1_ASAP7_75t_R%noxref_35
cc_243 N_noxref_35_1 N_MM24_g 0.00148871f
cc_244 N_noxref_35_1 N_QN_7 0.0383057f
x_PM_SDFLx1_ASAP7_75t_R%PD5 VSS N_MM17_s N_MM16_d N_PD5_1 N_PD5_4 N_PD5_5
+ PM_SDFLx1_ASAP7_75t_R%PD5
cc_245 N_PD5_1 N_MM18_g 0.000800328f
cc_246 N_PD5_4 N_MM18_g 0.00695307f
cc_247 N_PD5_5 N_MM18_g 0.0239955f
cc_248 N_PD5_4 N_MM17_g 0.0152564f
cc_249 N_PD5_1 N_MM16_g 0.000917171f
cc_250 N_PD5_5 N_MM16_g 0.0155834f
cc_251 N_PD5_1 N_SH_13 0.000513755f
cc_252 N_PD5_1 N_SH_15 0.000503119f
cc_253 N_PD5_1 N_SH_16 0.000570214f
cc_254 N_PD5_4 N_SH_5 0.000659341f
cc_255 N_PD5_1 N_SH_22 0.00240217f
x_PM_SDFLx1_ASAP7_75t_R%QN VSS QN N_MM24_d N_MM25_d N_QN_10 N_QN_7 N_QN_11
+ N_QN_2 N_QN_1 N_QN_8 N_QN_9 PM_SDFLx1_ASAP7_75t_R%QN
cc_256 N_QN_10 N_MM0_g 6.71559e-20
cc_257 N_QN_10 N_SE_9 0.000730087f
cc_258 N_QN_10 N_SE_13 0.000245287f
cc_259 N_QN_10 N_SE_12 0.00160811f
cc_260 N_QN_7 N_SH_20 0.00133324f
cc_261 N_QN_11 N_SH_25 0.000727563f
cc_262 N_QN_2 N_SH_2 0.000773655f
cc_263 N_QN_1 N_MM24_g 0.00120032f
cc_264 N_QN_2 N_MM24_g 0.00137805f
cc_265 N_QN_8 N_SH_2 0.001785f
cc_266 N_QN_8 N_MM24_g 0.0154711f
cc_267 N_QN_9 N_SH_20 0.00671346f
cc_268 N_QN_7 N_MM24_g 0.054339f
x_PM_SDFLx1_ASAP7_75t_R%noxref_36 VSS N_noxref_36_1
+ PM_SDFLx1_ASAP7_75t_R%noxref_36
cc_269 N_noxref_36_1 N_MM24_g 0.00149235f
cc_270 N_noxref_36_1 N_QN_8 0.0385706f
cc_271 N_noxref_36_1 N_noxref_35_1 0.00177166f
x_PM_SDFLx1_ASAP7_75t_R%SEN VSS N_MM27_g N_MM0_d N_MM2_d N_SEN_3 N_SEN_4
+ N_SEN_13 N_SEN_14 N_SEN_1 N_SEN_15 N_SEN_11 N_SEN_12 N_SEN_10 N_SEN_16
+ PM_SDFLx1_ASAP7_75t_R%SEN
cc_272 N_SEN_3 N_SE_9 0.000160716f
cc_273 N_SEN_4 N_SE_9 0.000174094f
cc_274 N_SEN_13 N_SE_9 0.00806088f
cc_275 N_SEN_14 N_SE_13 0.000228547f
cc_276 N_SEN_1 N_SE_8 0.000351449f
cc_277 N_SEN_15 N_SE_9 0.000407098f
cc_278 N_SEN_13 N_SE_12 0.000437889f
cc_279 N_SEN_11 N_MM0_g 0.0157398f
cc_280 N_SEN_12 N_SE_13 0.000464382f
cc_281 N_SEN_10 N_MM0_g 0.0537429f
cc_282 N_SEN_1 N_SE_1 0.00130748f
cc_283 N_SEN_13 N_SE_13 0.000517868f
cc_284 N_SEN_4 N_SE_2 0.000672221f
cc_285 N_SEN_4 N_MM0_g 0.00134222f
cc_286 N_SEN_12 N_SE_8 0.00174139f
cc_287 N_SEN_3 N_MM0_g 0.00175125f
cc_288 N_SEN_11 N_SE_2 0.00187685f
cc_289 N_MM27_g N_MM31_g 0.00330746f
cc_290 N_SEN_16 N_SE_13 0.0632777f
x_PM_SDFLx1_ASAP7_75t_R%SS VSS N_MM16_g N_MM14_d N_MM15_d N_SS_13 N_SS_15
+ N_SS_14 N_SS_17 N_SS_16 N_SS_12 N_SS_3 N_SS_4 N_SS_1 N_SS_11 N_SS_10
+ PM_SDFLx1_ASAP7_75t_R%SS
cc_291 N_MM16_g N_CLKN_10 0.000646394f
cc_292 N_MM16_g N_CLKN_5 0.000428827f
cc_293 N_MM16_g N_MM18_g 0.0133574f
cc_294 N_SS_13 N_SE_13 0.000911835f
cc_295 N_SS_15 N_SE_13 0.00320116f
cc_296 N_SS_14 N_SEN_3 0.00158983f
cc_297 N_SS_14 N_SEN_11 0.000114456f
cc_298 N_SS_14 N_SEN_15 0.000122262f
cc_299 N_SS_14 N_SEN_4 0.000266664f
cc_300 N_SS_13 N_SEN_16 0.000361669f
cc_301 N_SS_17 N_SEN_13 0.000379985f
cc_302 N_SS_16 N_SEN_15 0.000836078f
cc_303 N_SS_12 N_SEN_16 0.00251717f
cc_304 N_SS_14 N_SEN_13 0.00863272f
x_PM_SDFLx1_ASAP7_75t_R%MS VSS N_MM11_g N_MM6_d N_MM12_d N_MM7_d N_MM13_d
+ N_MS_3 N_MS_15 N_MS_12 N_MS_13 N_MS_1 N_MS_17 N_MS_4 N_MS_11 N_MS_18 N_MS_19
+ N_MS_14 N_MS_16 PM_SDFLx1_ASAP7_75t_R%MS
cc_305 N_MS_3 N_MM18_g 5.88759e-20
cc_306 N_MS_3 N_CLKN_29 0.00015076f
cc_307 N_MS_3 N_CLKN_10 0.000657117f
cc_308 N_MS_3 N_CLKN_3 9.2419e-20
cc_309 N_MS_3 N_CLKN_35 0.000138297f
cc_310 N_MS_15 N_CLKN_29 0.000280515f
cc_311 N_MS_12 N_MM12_g 0.00787602f
cc_312 N_MS_13 N_MM12_g 0.00779411f
cc_313 N_MS_15 N_CLKN_10 0.000386934f
cc_314 N_MS_1 N_MM9_g 0.000692827f
cc_315 N_MS_17 N_CLKN_10 0.00158737f
cc_316 N_MS_4 N_MM12_g 0.00230808f
cc_317 N_MS_11 N_MM12_g 0.00651622f
cc_318 N_MS_4 N_CLKN_10 0.00638196f
cc_319 N_MM11_g N_MM9_g 0.0141603f
cc_320 N_MS_3 N_MM12_g 0.0259458f
cc_321 N_MS_18 N_SEN_16 0.000868003f
cc_322 N_MS_19 N_SEN_16 0.00298721f
cc_323 N_MS_13 N_CLKB_22 0.00035323f
cc_324 N_MS_13 N_MM10_g 0.000138152f
cc_325 N_MS_13 N_CLKB_18 0.00017752f
cc_326 N_MS_13 N_CLKB_2 0.00019557f
cc_327 N_MS_17 N_CLKB_18 0.00422954f
cc_328 N_MS_17 N_CLKB_2 0.00037142f
cc_329 N_MS_19 N_CLKB_18 0.00040803f
cc_330 N_MS_18 N_CLKB_22 0.00160484f
cc_331 N_MS_13 N_MM17_g 0.0154329f
x_PM_SDFLx1_ASAP7_75t_R%SE VSS SE N_MM31_g N_MM0_g N_SE_9 N_SE_13 N_SE_8
+ N_SE_12 N_SE_1 N_SE_2 N_SE_10 N_SE_7 N_SE_11 PM_SDFLx1_ASAP7_75t_R%SE
x_PM_SDFLx1_ASAP7_75t_R%SH VSS N_MM14_g N_MM24_g N_MM13_s N_MM18_d N_MM12_s
+ N_MM17_d N_SH_14 N_SH_25 N_SH_21 N_SH_23 N_SH_6 N_SH_13 N_SH_18 N_SH_16
+ N_SH_17 N_SH_5 N_SH_22 N_SH_20 N_SH_2 N_SH_15 N_SH_1 N_SH_19 N_SH_24
+ PM_SDFLx1_ASAP7_75t_R%SH
cc_332 N_SH_14 N_CLKN_35 9.17988e-20
cc_333 N_SH_25 N_CLKN_10 9.21541e-20
cc_334 N_SH_21 N_CLKN_10 0.000199637f
cc_335 N_SH_23 N_CLKN_10 0.000212381f
cc_336 N_SH_6 N_CLKN_10 0.000256826f
cc_337 N_SH_13 N_MM12_g 0.00677829f
cc_338 N_SH_18 N_CLKN_10 0.000388114f
cc_339 N_SH_16 N_CLKN_10 0.000446605f
cc_340 N_SH_17 N_CLKN_10 0.000564633f
cc_341 N_SH_14 N_CLKN_5 0.000674955f
cc_342 N_SH_6 N_MM18_g 0.00100479f
cc_343 N_SH_5 N_CLKN_10 0.00283521f
cc_344 N_SH_5 N_MM12_g 0.00948043f
cc_345 N_SH_14 N_MM18_g 0.0161929f
cc_346 N_SH_22 N_SE_13 0.000221105f
cc_347 N_SH_20 N_SE_12 0.000226514f
cc_348 N_SH_2 N_SE_2 0.0016708f
cc_349 N_SH_15 N_SE_13 0.00103025f
cc_350 N_SH_25 N_SE_13 0.00215637f
cc_351 N_SH_16 N_SE_13 0.00271258f
cc_352 N_MM24_g N_MM0_g 0.00331022f
cc_353 N_SH_20 N_SE_9 0.00577647f
cc_354 N_SH_1 N_SEN_3 0.000213211f
cc_355 N_MM24_g N_SEN_4 9.91647e-20
cc_356 N_SH_25 N_SEN_15 0.000106923f
cc_357 N_MM14_g N_SEN_3 0.000113303f
cc_358 N_SH_20 N_SEN_4 0.000161138f
cc_359 N_SH_25 N_SEN_13 0.00150765f
cc_360 N_SH_18 N_SEN_16 0.000180979f
cc_361 N_MM24_g N_SEN_3 0.00019343f
cc_362 N_SH_20 N_SEN_15 0.000255779f
cc_363 N_SH_19 N_SEN_16 0.000321248f
cc_364 N_SH_15 N_SEN_16 0.000377016f
cc_365 N_SH_25 N_SEN_16 0.00481277f
cc_366 N_SH_16 N_SEN_16 0.00604355f
cc_367 N_SH_6 N_MM17_g 0.000164949f
cc_368 N_SH_14 N_MM17_g 0.00675461f
cc_369 N_SH_13 N_MM17_g 0.00679153f
cc_370 N_SH_21 N_CLKB_18 0.000294438f
cc_371 N_SH_15 N_CLKB_18 0.000381738f
cc_372 N_SH_17 N_CLKB_18 0.000450062f
cc_373 N_SH_16 N_CLKB_2 0.000478169f
cc_374 N_SH_5 N_CLKB_2 0.000500678f
cc_375 N_SH_23 N_CLKB_18 0.000503205f
cc_376 N_SH_25 N_CLKB_22 0.000899228f
cc_377 N_SH_16 N_CLKB_18 0.00453078f
cc_378 N_SH_15 N_CLKB_22 0.00107025f
cc_379 N_SH_5 N_MM17_g 0.0183709f
cc_380 N_SH_17 N_MS_3 9.9312e-20
cc_381 N_SH_21 N_MS_3 0.000181673f
cc_382 N_SH_6 N_MS_3 0.00021626f
cc_383 N_SH_14 N_MS_3 0.000436505f
cc_384 N_SH_13 N_MS_3 0.000231694f
cc_385 N_SH_13 N_MS_11 0.000233146f
cc_386 N_SH_21 N_MS_4 0.000313578f
cc_387 N_SH_15 N_MS_16 0.000405471f
cc_388 N_SH_6 N_MS_4 0.000417682f
cc_389 N_SH_21 N_MS_17 0.000537518f
cc_390 N_SH_14 N_MS_4 0.000608238f
cc_391 N_SH_15 N_MS_19 0.00133351f
cc_392 N_SH_5 N_MS_3 0.00371277f
cc_393 N_SH_17 N_MM16_g 0.000104471f
cc_394 N_SH_19 N_MM16_g 0.000311383f
cc_395 N_MM14_g N_SS_3 0.000315775f
cc_396 N_MM14_g N_SS_4 0.000420905f
cc_397 N_SH_22 N_SS_15 0.000584084f
cc_398 N_SH_24 N_SS_16 0.000663004f
cc_399 N_SH_24 N_SS_14 0.000807854f
cc_400 N_SH_16 N_SS_1 0.00081088f
cc_401 N_SH_1 N_SS_14 0.000884895f
cc_402 N_MM14_g N_SS_1 0.0011143f
cc_403 N_SH_1 N_MM16_g 0.00129795f
cc_404 N_SH_18 N_SS_12 0.00149463f
cc_405 N_SH_25 N_SS_14 0.00178257f
cc_406 N_MM14_g N_SS_11 0.00655832f
cc_407 N_MM14_g N_SS_10 0.00659453f
cc_408 N_SH_16 N_SS_12 0.00446197f
cc_409 N_SH_19 N_SS_14 0.00482636f
cc_410 N_MM14_g N_MM16_g 0.0299881f
x_PM_SDFLx1_ASAP7_75t_R%CLKB VSS N_MM10_g N_MM17_g N_MM23_d N_MM22_d N_CLKB_13
+ N_CLKB_22 N_CLKB_16 N_CLKB_5 N_CLKB_19 N_CLKB_15 N_CLKB_6 N_CLKB_20 N_CLKB_14
+ N_CLKB_17 N_CLKB_18 N_CLKB_2 N_CLKB_1 N_CLKB_21 PM_SDFLx1_ASAP7_75t_R%CLKB
cc_411 N_CLKB_13 N_CLK_5 7.96528e-20
cc_412 N_CLKB_22 N_CLK_5 0.000113309f
cc_413 N_CLKB_16 N_CLK_5 0.000539518f
cc_414 N_CLKB_5 N_CLK_5 0.00036059f
cc_415 N_CLKB_19 N_CLK_5 0.00220891f
cc_416 N_CLKB_22 N_CLKN_10 2.72031e-20
cc_417 N_CLKB_22 N_CLKN_8 3.20588e-20
cc_418 N_CLKB_22 N_CLKN_25 3.2796e-20
cc_419 N_CLKB_22 N_MM22_g 4.88099e-20
cc_420 N_CLKB_5 N_CLKN_23 7.9392e-20
cc_421 N_CLKB_15 N_CLKN_26 9.30476e-20
cc_422 N_CLKB_19 N_CLKN_27 0.000109984f
cc_423 N_CLKB_6 N_CLKN_33 0.000172854f
cc_424 N_MM17_g N_CLKN_5 0.000199228f
cc_425 N_CLKB_20 N_CLKN_33 0.000258416f
cc_426 N_CLKB_22 N_CLKN_29 0.000659916f
cc_427 N_CLKB_22 N_CLKN_28 0.000328036f
cc_428 N_CLKB_14 N_MM22_g 0.0112188f
cc_429 N_CLKB_13 N_MM22_g 0.0385771f
cc_430 N_CLKB_15 N_CLKN_27 0.000366651f
cc_431 N_CLKB_17 N_CLKN_35 0.000478463f
cc_432 N_CLKB_18 N_CLKN_10 0.000524093f
cc_433 N_MM10_g N_CLKN_3 0.000559239f
cc_434 N_CLKB_5 N_MM22_g 0.000584722f
cc_435 N_CLKB_16 N_CLKN_1 0.000589463f
cc_436 N_CLKB_16 N_CLKN_35 0.000620606f
cc_437 N_CLKB_2 N_CLKN_10 0.00269591f
cc_438 N_CLKB_1 N_CLKN_2 0.00214545f
cc_439 N_CLKB_14 N_CLKN_1 0.000838963f
cc_440 N_CLKB_6 N_MM22_g 0.000848157f
cc_441 N_MM10_g N_MM1_g 0.00164299f
cc_442 N_CLKB_21 N_CLKN_34 0.00181744f
cc_443 N_CLKB_17 N_CLKN_28 0.00263077f
cc_444 N_CLKB_15 N_CLKN_33 0.00354991f
cc_445 N_CLKB_16 N_CLKN_27 0.00472052f
cc_446 N_MM17_g N_CLKN_10 0.00496732f
cc_447 N_MM17_g N_MM12_g 0.00566544f
cc_448 N_MM10_g N_MM9_g 0.00909902f
cc_449 N_MM17_g N_MM18_g 0.0184151f
cc_450 N_CLKB_22 N_CLKN_35 0.0458367f
cc_451 N_CLKB_16 N_SE_1 5.78543e-20
cc_452 N_CLKB_5 N_SE_10 5.90055e-20
cc_453 N_CLKB_5 N_SE_7 0.000179503f
cc_454 N_CLKB_16 N_SE_7 0.0033304f
cc_455 N_CLKB_18 N_SE_13 0.000495508f
cc_456 N_CLKB_19 N_SE_10 0.00174478f
cc_457 N_CLKB_22 N_SE_13 0.00234408f
cc_458 N_CLKB_22 N_SE_8 0.00361589f
cc_459 N_CLKB_16 N_SE_11 0.0063228f
cc_460 N_CLKB_22 N_SEN_12 0.00408441f
cc_461 N_CLKB_18 N_SEN_16 0.00291908f
cc_462 N_CLKB_17 N_SEN_16 0.000336414f
cc_463 N_CLKB_22 N_SEN_16 0.00996458f
cc_464 N_CLKB_22 N_SI_4 0.00249093f
x_PM_SDFLx1_ASAP7_75t_R%CLKN VSS N_MM22_g N_MM1_g N_MM9_g N_MM12_g N_MM18_g
+ N_MM20_d N_MM21_d N_CLKN_30 N_CLKN_27 N_CLKN_26 N_CLKN_31 N_CLKN_8 N_CLKN_33
+ N_CLKN_21 N_CLKN_22 N_CLKN_1 N_CLKN_9 N_CLKN_35 N_CLKN_25 N_CLKN_23 N_CLKN_2
+ N_CLKN_28 N_CLKN_34 N_CLKN_10 N_CLKN_5 N_CLKN_29 N_CLKN_3 N_CLKN_32 N_CLKN_24
+ PM_SDFLx1_ASAP7_75t_R%CLKN
cc_465 N_CLKN_30 N_MM20_g 6.89415e-20
cc_466 N_CLKN_27 N_MM20_g 6.93672e-20
cc_467 N_CLKN_26 N_MM20_g 8.89276e-20
cc_468 N_CLKN_31 N_MM20_g 9.79398e-20
cc_469 N_CLKN_8 N_MM20_g 0.00112459f
cc_470 N_CLKN_33 N_MM20_g 0.00034696f
cc_471 N_CLKN_21 N_MM20_g 0.0112099f
cc_472 N_CLKN_22 N_MM20_g 0.0113154f
cc_473 N_CLKN_31 N_CLK_4 0.000405093f
cc_474 N_CLKN_1 N_CLK_6 0.0005874f
cc_475 N_CLKN_9 N_MM20_g 0.000640698f
cc_476 N_CLKN_35 N_CLK_4 0.000670927f
cc_477 N_CLKN_27 N_CLK_6 0.000944507f
cc_478 N_CLKN_25 N_CLK_6 0.000954175f
cc_479 N_CLKN_1 N_CLK_1 0.0035354f
cc_480 N_CLKN_23 N_CLK_4 0.00165569f
cc_481 N_CLKN_25 N_CLK_5 0.00169422f
cc_482 N_CLKN_27 N_CLK_4 0.00461393f
cc_483 N_MM22_g N_MM20_g 0.0350789f
*END of SDFLx1_ASAP7_75t_R.pxi
.ENDS
** Design:	SDFLx2_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "SDFLx2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "SDFLx2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_SDFLx2_ASAP7_75t_R%NET0168 VSS 2 3 1
c1 1 VSS 0.000995471f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3780 $Y2=0.0675
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%noxref_34 VSS 1
c1 1 VSS 0.00477386f
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%noxref_33 VSS 1
c1 1 VSS 0.00446376f
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%D VSS 4 3 1 5
c1 1 VSS 0.00723928f
c2 3 VSS 0.0462111f
c3 4 VSS 0.00464072f
c4 5 VSS 0.00368478f
r1 5 7 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.1080 $X2=0.4050 $Y2=0.1215
r2 4 7 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1215
r3 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r4 4 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%PD3 VSS 2 4 1
c1 1 VSS 0.00091033f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.0405 $X2=0.7065 $Y2=0.0405
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.0405 $X2=0.6895 $Y2=0.0405
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6895 $Y=0.0405 $X2=0.7065 $Y2=0.0405
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%PD4 VSS 2 4 1
c1 1 VSS 0.00102999f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9890 $Y=0.2295 $X2=0.9765 $Y2=0.2295
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9550 $Y=0.2295 $X2=0.9595 $Y2=0.2295
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9595 $Y=0.2295 $X2=0.9765 $Y2=0.2295
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%NET0144 VSS 12 13 27 28 9 7 1 2 8
c1 1 VSS 0.00533332f
c2 2 VSS 0.00531469f
c3 7 VSS 0.0033348f
c4 8 VSS 0.00335745f
c5 9 VSS 0.00273696f
r1 28 26 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r2 2 26 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r4 27 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r5 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4280 $Y2=0.1980
r6 21 22 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4185
+ $Y=0.1980 $X2=0.4280 $Y2=0.1980
r7 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1980 $X2=0.4185 $Y2=0.1980
r8 19 20 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.3875
+ $Y=0.1980 $X2=0.4050 $Y2=0.1980
r9 18 19 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3695
+ $Y=0.1980 $X2=0.3875 $Y2=0.1980
r10 17 18 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1980 $X2=0.3695 $Y2=0.1980
r11 16 17 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.1980 $X2=0.3510 $Y2=0.1980
r12 15 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1980 $X2=0.3375 $Y2=0.1980
r13 14 15 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3130
+ $Y=0.1980 $X2=0.3240 $Y2=0.1980
r14 9 14 0.699569 $w=1.3e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.3100
+ $Y=0.1980 $X2=0.3130 $Y2=0.1980
r15 1 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.1980
r16 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r17 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r18 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r19 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.00423273f
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.00424703f
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%PU1 VSS 13 24 26 10 2 11 8 1 9
c1 1 VSS 0.00650247f
c2 2 VSS 0.00859773f
c3 8 VSS 0.00354247f
c4 9 VSS 0.00237496f
c5 10 VSS 0.00216341f
c6 11 VSS 0.0231065f
r1 26 25 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r2 10 25 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5420 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r3 9 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4840 $Y2=0.2025
r4 24 9 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r5 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5130 $Y=0.2025
+ $X2=0.4900 $Y2=0.2340
r6 20 21 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4810
+ $Y=0.2340 $X2=0.4900 $Y2=0.2340
r7 19 20 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4690
+ $Y=0.2340 $X2=0.4810 $Y2=0.2340
r8 18 19 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4540
+ $Y=0.2340 $X2=0.4690 $Y2=0.2340
r9 17 18 17.7224 $w=1.3e-08 $l=7.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.4540 $Y2=0.2340
r10 16 17 19.5879 $w=1.3e-08 $l=8.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2940
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r11 15 16 5.59655 $w=1.3e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.2940 $Y2=0.2340
r12 11 15 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2580
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r13 8 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2160
+ $X2=0.2700 $Y2=0.2340
r14 1 8 23.8708 $w=2.02e-08 $l=4.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.2700 $Y=0.1755 $X2=0.2700 $Y2=0.2160
r15 13 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r16 8 12 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r17 2 10 1e-05
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%CLK VSS 11 3 4 6 1 5
c1 1 VSS 0.00307103f
c2 3 VSS 0.0599236f
c3 4 VSS 0.00149615f
c4 5 VSS 0.00465296f
c5 6 VSS 0.0019696f
r1 5 14 4.60559 $w=1.39091e-08 $l=2.74591e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0630 $X2=0.1030 $Y2=0.0900
r2 13 14 1.45753 $w=1.53529e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.0900 $X2=0.1030 $Y2=0.0900
r3 6 13 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0900 $X2=0.0945 $Y2=0.0900
r4 11 10 0.757867 $w=1.3e-08 $l=3.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1500 $X2=0.0810 $Y2=0.1467
r5 9 10 2.73998 $w=1.3e-08 $l=1.17e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1467
r6 8 9 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1235 $X2=0.0810 $Y2=0.1350
r7 4 8 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1100 $X2=0.0810 $Y2=0.1235
r8 4 6 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1100 $X2=0.0810 $Y2=0.0900
r9 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r10 1 9 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%noxref_29 VSS 1
c1 1 VSS 0.00582343f
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%noxref_27 VSS 1
c1 1 VSS 0.00437018f
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%PD2 VSS 7 12 4 5 1
c1 1 VSS 0.00742609f
c2 4 VSS 0.00184285f
c3 5 VSS 0.00234061f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7040 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r3 9 5 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.6765
+ $Y=0.2295 $X2=0.7020 $Y2=0.2295
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.6615
+ $Y=0.2295 $X2=0.6765 $Y2=0.2295
r5 1 8 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.6480
+ $Y=0.2295 $X2=0.6615 $Y2=0.2295
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.2295 $X2=0.6460 $Y2=0.2295
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.2295 $X2=0.6335 $Y2=0.2295
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%noxref_35 VSS 1
c1 1 VSS 0.0423952f
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%noxref_32 VSS 1
c1 1 VSS 0.00370373f
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%noxref_31 VSS 1
c1 1 VSS 0.00347143f
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%SS VSS 9 34 39 13 15 14 17 16 12 3 4 1 10 11
c1 1 VSS 0.0011126f
c2 3 VSS 0.00556991f
c3 4 VSS 0.0066391f
c4 9 VSS 0.0384173f
c5 10 VSS 0.00349756f
c6 11 VSS 0.00365109f
c7 12 VSS 0.000996111f
c8 13 VSS 0.00845762f
c9 14 VSS 0.00177281f
c10 15 VSS 0.00251824f
c11 16 VSS 0.00603784f
c12 17 VSS 0.00224605f
r1 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0655 $Y=0.2295 $X2=1.0780 $Y2=0.2295
r2 39 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0630 $Y=0.2295 $X2=1.0655 $Y2=0.2295
r3 4 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0800 $Y=0.2295
+ $X2=1.0800 $Y2=0.2340
r4 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.0800
+ $Y=0.2340 $X2=1.0935 $Y2=0.2340
r5 16 32 7.21452 $w=1.425e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.2340 $X2=1.1070 $Y2=0.1980
r6 16 37 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1070 $Y=0.2340 $X2=1.0935 $Y2=0.2340
r7 10 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.0655 $Y=0.0405 $X2=1.0780 $Y2=0.0405
r8 34 10 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.0630 $Y=0.0405 $X2=1.0655 $Y2=0.0405
r9 31 32 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.1440 $X2=1.1070 $Y2=0.1980
r10 14 30 8.95608 $w=1.36627e-08 $l=4.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1070 $Y=0.0810 $X2=1.1070 $Y2=0.0395
r11 14 31 14.691 $w=1.3e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.0810 $X2=1.1070 $Y2=0.1440
r12 3 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0800 $Y=0.0405
+ $X2=1.0800 $Y2=0.0360
r13 17 29 1.40651 $w=1.51875e-08 $l=1.45774e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1070 $Y=0.0305 $X2=1.0935 $Y2=0.0360
r14 17 30 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.0305 $X2=1.1070 $Y2=0.0395
r15 28 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.0800
+ $Y=0.0360 $X2=1.0935 $Y2=0.0360
r16 27 28 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.0685
+ $Y=0.0360 $X2=1.0800 $Y2=0.0360
r17 26 27 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.0640
+ $Y=0.0360 $X2=1.0685 $Y2=0.0360
r18 25 26 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.0360 $X2=1.0640 $Y2=0.0360
r19 13 15 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0260 $Y=0.0360 $X2=0.9990 $Y2=0.0360
r20 13 25 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.0360 $X2=1.0530 $Y2=0.0360
r21 12 22 8.04505 $w=1.3e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.9990
+ $Y=0.0705 $X2=0.9990 $Y2=0.1050
r22 12 15 6.39593 $w=1.55565e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9990 $Y=0.0705 $X2=0.9990 $Y2=0.0360
r23 1 19 2.36633 $w=2.3e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.9990
+ $Y=0.1055 $X2=0.9990 $Y2=0.1055
r24 1 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.9990 $Y=0.1055
+ $X2=0.9990 $Y2=0.1050
r25 9 19 0.314665 $w=2.27e-07 $l=2.95e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.9990 $Y=0.1350 $X2=0.9990 $Y2=0.1055
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%noxref_36 VSS 1
c1 1 VSS 0.0423525f
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%PD5 VSS 7 12 1 5 4
c1 1 VSS 0.00743021f
c2 4 VSS 0.00187932f
c3 5 VSS 0.00237028f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9890 $Y=0.0405 $X2=0.9865 $Y2=0.0405
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9740 $Y=0.0405 $X2=0.9865 $Y2=0.0405
r3 9 5 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.9585
+ $Y=0.0405 $X2=0.9720 $Y2=0.0405
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.9435
+ $Y=0.0405 $X2=0.9585 $Y2=0.0405
r5 1 8 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.9180
+ $Y=0.0405 $X2=0.9435 $Y2=0.0405
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9035 $Y=0.0405 $X2=0.9160 $Y2=0.0405
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9010 $Y=0.0405 $X2=0.9035 $Y2=0.0405
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%QN VSS 22 16 17 28 29 9 7 8 10 11 1 2
c1 1 VSS 0.0101587f
c2 2 VSS 0.0104033f
c3 7 VSS 0.0045053f
c4 8 VSS 0.00449869f
c5 9 VSS 0.00922717f
c6 10 VSS 0.00918285f
c7 11 VSS 0.00729022f
c8 12 VSS 0.00338348f
c9 13 VSS 0.00334621f
r1 29 27 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.3130 $Y=0.2025 $X2=1.3105 $Y2=0.2025
r2 2 27 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.2960 $Y=0.2025 $X2=1.3105 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.2815 $Y=0.2025 $X2=1.2960 $Y2=0.2025
r4 28 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.2790 $Y=0.2025 $X2=1.2815 $Y2=0.2025
r5 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.2960 $Y=0.2025
+ $X2=1.2960 $Y2=0.2340
r6 24 25 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=1.2960
+ $Y=0.2340 $X2=1.3365 $Y2=0.2340
r7 10 24 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.2845
+ $Y=0.2340 $X2=1.2960 $Y2=0.2340
r8 13 23 0.624487 $w=2.20462e-08 $l=9.8e-09 $layer=M1 $thickness=3.6e-08
+ $X=1.3770 $Y=0.2340 $X2=1.3770 $Y2=0.2242
r9 13 25 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3770 $Y=0.2340 $X2=1.3365 $Y2=0.2340
r10 22 23 0.291487 $w=1.3e-08 $l=1.2e-09 $layer=M1 $thickness=3.6e-08 $X=1.3770
+ $Y=0.2230 $X2=1.3770 $Y2=0.2242
r11 22 21 2.73998 $w=1.3e-08 $l=1.18e-08 $layer=M1 $thickness=3.6e-08 $X=1.3770
+ $Y=0.2230 $X2=1.3770 $Y2=0.2112
r12 20 21 15.4488 $w=1.3e-08 $l=6.62e-08 $layer=M1 $thickness=3.6e-08 $X=1.3770
+ $Y=0.1450 $X2=1.3770 $Y2=0.2112
r13 11 12 5.69636 $w=1.58e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3770 $Y=0.0675 $X2=1.3770 $Y2=0.0360
r14 11 20 18.0722 $w=1.3e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=1.3770
+ $Y=0.0675 $X2=1.3770 $Y2=0.1450
r15 12 19 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3770 $Y=0.0360 $X2=1.3365 $Y2=0.0360
r16 18 19 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=1.2960
+ $Y=0.0360 $X2=1.3365 $Y2=0.0360
r17 9 18 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.2845
+ $Y=0.0360 $X2=1.2960 $Y2=0.0360
r18 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.2960 $Y=0.0675
+ $X2=1.2960 $Y2=0.0360
r19 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.3130 $Y=0.0675 $X2=1.3105 $Y2=0.0675
r20 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.2960 $Y=0.0675 $X2=1.3105 $Y2=0.0675
r21 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.2815 $Y=0.0675 $X2=1.2960 $Y2=0.0675
r22 16 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.2790 $Y=0.0675 $X2=1.2815 $Y2=0.0675
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%MH VSS 9 55 59 62 66 10 3 21 17 1 4 12 14 18 20
+ 16 19 15
c1 1 VSS 0.000217514f
c2 3 VSS 0.00473607f
c3 4 VSS 0.00495982f
c4 9 VSS 0.0361308f
c5 10 VSS 0.00227007f
c6 11 VSS 9.98988e-20
c7 12 VSS 0.00211122f
c8 13 VSS 6.71813e-20
c9 14 VSS 0.00937465f
c10 15 VSS 0.00780178f
c11 16 VSS 0.00174677f
c12 17 VSS 0.00061796f
c13 18 VSS 0.000936186f
c14 19 VSS 0.00298503f
c15 20 VSS 5.93629e-20
c16 21 VSS 0.00269034f
r1 66 65 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.2295 $X2=0.6085 $Y2=0.2295
r2 64 65 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6040 $Y=0.2295 $X2=0.6085 $Y2=0.2295
r3 3 64 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5920 $Y=0.2295 $X2=0.6040 $Y2=0.2295
r4 13 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2295 $X2=0.5920 $Y2=0.2295
r5 60 61 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.1890 $X2=0.5840 $Y2=0.1890
r6 62 60 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.1890 $X2=0.5795 $Y2=0.1890
r7 12 61 0.185185 $w=5.4e-08 $l=1e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.1890 $X2=0.5840 $Y2=0.1890
r8 12 3 0.518519 $w=3.9e-08 $l=4.05494e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.1890 $X2=0.5920 $Y2=0.2295
r9 59 58 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r10 57 58 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6580 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r11 4 57 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6460 $Y=0.0405 $X2=0.6580 $Y2=0.0405
r12 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0405 $X2=0.6460 $Y2=0.0405
r13 10 4 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0810 $X2=0.6460 $Y2=0.0810
r14 55 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.0810 $X2=0.6335 $Y2=0.0810
r15 3 47 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2295
+ $X2=0.5900 $Y2=0.2340
r16 4 41 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.0405
+ $X2=0.6440 $Y2=0.0360
r17 44 45 1.63233 $w=1.3e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.5990
+ $Y=0.2340 $X2=0.6060 $Y2=0.2340
r18 44 47 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5990
+ $Y=0.2340 $X2=0.5900 $Y2=0.2340
r19 43 45 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.6105
+ $Y=0.2340 $X2=0.6060 $Y2=0.2340
r20 42 43 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6305
+ $Y=0.2340 $X2=0.6105 $Y2=0.2340
r21 14 21 4.53042 $w=1.46981e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6665 $Y=0.2340 $X2=0.6930 $Y2=0.2340
r22 14 42 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.6665
+ $Y=0.2340 $X2=0.6305 $Y2=0.2340
r23 15 39 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.6530
+ $Y=0.0360 $X2=0.6705 $Y2=0.0360
r24 15 41 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6530
+ $Y=0.0360 $X2=0.6440 $Y2=0.0360
r25 21 38 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.2340 $X2=0.6930 $Y2=0.2160
r26 19 33 2.43171 $w=1.804e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6930 $Y=0.0360 $X2=0.6930 $Y2=0.0535
r27 19 39 3.59766 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.0360 $X2=0.6705 $Y2=0.0360
r28 37 38 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1980 $X2=0.6930 $Y2=0.2160
r29 36 37 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1800 $X2=0.6930 $Y2=0.1980
r30 35 36 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1680 $X2=0.6930 $Y2=0.1800
r31 34 35 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1590 $X2=0.6930 $Y2=0.1680
r32 17 20 2.43413 $w=1.59032e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6930 $Y=0.1465 $X2=0.6930 $Y2=0.1310
r33 17 34 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1465 $X2=0.6930 $Y2=0.1590
r34 32 33 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.0625 $X2=0.6930 $Y2=0.0535
r35 31 32 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.0720 $X2=0.6930 $Y2=0.0625
r36 30 31 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.0900 $X2=0.6930 $Y2=0.0720
r37 29 30 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1025 $X2=0.6930 $Y2=0.0900
r38 16 20 2.78392 $w=1.56471e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6930 $Y=0.1140 $X2=0.6930 $Y2=0.1310
r39 16 29 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1140 $X2=0.6930 $Y2=0.1025
r40 20 28 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1310 $X2=0.7110 $Y2=0.1310
r41 27 28 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1310 $X2=0.7110 $Y2=0.1310
r42 18 26 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.1310 $X2=0.7830 $Y2=0.1310
r43 18 27 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.1310 $X2=0.7290 $Y2=0.1310
r44 1 23 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.7830
+ $Y=0.1310 $X2=0.7830 $Y2=0.1310
r45 1 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7830 $Y=0.1310
+ $X2=0.7830 $Y2=0.1310
r46 9 23 0.314665 $w=2.27e-07 $l=4e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.7830 $Y=0.1350 $X2=0.7830 $Y2=0.1310
r47 3 12 1e-05
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%MS VSS 10 43 46 50 52 3 15 13 12 1 17 11 4 18 19
+ 14 16
c1 1 VSS 0.00317613f
c2 3 VSS 0.00575041f
c3 4 VSS 0.00955867f
c4 10 VSS 0.0376965f
c5 11 VSS 0.00331324f
c6 12 VSS 0.00314415f
c7 13 VSS 0.00265374f
c8 14 VSS 0.000855988f
c9 15 VSS 0.00355279f
c10 16 VSS 0.00188635f
c11 17 VSS 0.00113231f
c12 18 VSS 0.00137182f
c13 19 VSS 0.00118316f
c14 20 VSS 0.00294966f
r1 52 51 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8810 $Y=0.2295 $X2=0.8785 $Y2=0.2295
r2 13 51 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8660 $Y=0.2295 $X2=0.8785 $Y2=0.2295
r3 12 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.2295 $X2=0.8080 $Y2=0.2295
r4 50 12 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.2295 $X2=0.7955 $Y2=0.2295
r5 47 13 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8370 $Y=0.2295 $X2=0.8640 $Y2=0.2295
r6 4 47 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08 $X=0.8100
+ $Y=0.2295 $X2=0.8370 $Y2=0.2295
r7 4 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8100 $Y=0.2295
+ $X2=0.8100 $Y2=0.2340
r8 15 20 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.2340 $X2=0.8370 $Y2=0.2340
r9 46 45 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8270 $Y=0.0405 $X2=0.8245 $Y2=0.0405
r10 44 45 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8200 $Y=0.0405 $X2=0.8245 $Y2=0.0405
r11 3 44 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8080 $Y=0.0405 $X2=0.8200 $Y2=0.0405
r12 11 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.0405 $X2=0.8080 $Y2=0.0405
r13 43 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.0405 $X2=0.7955 $Y2=0.0405
r14 20 39 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.2340 $X2=0.8370 $Y2=0.2160
r15 3 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8100 $Y=0.0405
+ $X2=0.8100 $Y2=0.0535
r16 38 39 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1870 $X2=0.8370 $Y2=0.2160
r17 37 38 4.89699 $w=1.3e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1660 $X2=0.8370 $Y2=0.1870
r18 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1525 $X2=0.8370 $Y2=0.1660
r19 35 36 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1310 $X2=0.8370 $Y2=0.1525
r20 34 35 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1115 $X2=0.8370 $Y2=0.1310
r21 17 31 1.15159 $w=1.75e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1000 $X2=0.8370 $Y2=0.0900
r22 17 34 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1000 $X2=0.8370 $Y2=0.1115
r23 16 32 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0625 $X2=0.8100 $Y2=0.0720
r24 16 33 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0625 $X2=0.8100 $Y2=0.0535
r25 30 31 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8235 $Y=0.0900 $X2=0.8370 $Y2=0.0900
r26 19 28 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.0900 $X2=0.7965 $Y2=0.0900
r27 19 30 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.0900 $X2=0.8235 $Y2=0.0900
r28 19 32 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0900 $X2=0.8100 $Y2=0.0720
r29 27 28 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.7740
+ $Y=0.0900 $X2=0.7965 $Y2=0.0900
r30 14 27 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7470
+ $Y=0.0900 $X2=0.7740 $Y2=0.0900
r31 14 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7470 $Y=0.0900
+ $X2=0.7500 $Y2=0.0900
r32 14 18 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7470
+ $Y=0.0900 $X2=0.7290 $Y2=0.0900
r33 25 26 5.02115 $w=1.53e-08 $l=8.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.7415 $Y=0.0900 $X2=0.7500 $Y2=0.0900
r34 23 25 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.7385 $Y=0.0900 $X2=0.7415 $Y2=0.0900
r35 1 23 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.7285
+ $Y=0.0900 $X2=0.7385 $Y2=0.0900
r36 1 22 2.48102 $w=2.2e-08 $l=5e-10 $layer=LIG $thickness=4.8e-08 $X=0.7285
+ $Y=0.0900 $X2=0.7290 $Y2=0.0900
r37 22 25 1.47681 $w=1.53e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7290 $Y=0.0900 $X2=0.7415 $Y2=0.0900
r38 10 22 0.314665 $w=2.27e-07 $l=4.5e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.7290 $Y=0.1350 $X2=0.7290 $Y2=0.0900
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%CLKB VSS 11 12 61 63 13 22 16 5 19 15 6 20 14 17
+ 18 2 1 21
c1 1 VSS 0.00014784f
c2 2 VSS 0.000212919f
c3 5 VSS 0.00733834f
c4 6 VSS 0.00723995f
c5 11 VSS 0.00449171f
c6 12 VSS 0.00460296f
c7 13 VSS 0.00744581f
c8 14 VSS 0.00749568f
c9 15 VSS 0.00646136f
c10 16 VSS 0.00361238f
c11 17 VSS 0.000128199f
c12 18 VSS 0.000486522f
c13 19 VSS 0.00590523f
c14 20 VSS 0.0030599f
c15 21 VSS 0.000163927f
c16 22 VSS 0.0197171f
r1 14 6 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1600 $Y2=0.2160
r2 63 14 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r3 6 56 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r4 13 5 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1600 $Y2=0.0540
r5 61 13 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r6 56 57 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r7 15 56 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1505
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r8 5 53 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r9 20 49 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.1890 $Y2=0.2160
r10 20 57 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2340 $X2=0.1755 $Y2=0.2340
r11 53 54 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r12 19 44 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1890 $Y2=0.0630
r13 19 54 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1755 $Y2=0.0360
r14 1 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6210 $Y=0.1350
+ $X2=0.6210 $Y2=0.1395
r15 11 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1350
r16 48 49 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1980 $X2=0.1890 $Y2=0.2160
r17 47 48 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1765 $X2=0.1890 $Y2=0.1980
r18 46 47 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1630 $X2=0.1890 $Y2=0.1765
r19 45 46 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1530 $X2=0.1890 $Y2=0.1630
r20 43 44 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0900 $X2=0.1890 $Y2=0.0630
r21 42 43 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1100 $X2=0.1890 $Y2=0.0900
r22 16 42 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1325 $X2=0.1890 $Y2=0.1100
r23 16 45 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1325 $X2=0.1890 $Y2=0.1530
r24 21 39 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1620 $X2=0.6210 $Y2=0.1395
r25 21 33 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.6210 $Y=0.1620 $X2=0.6210
+ $Y2=0.1530
r26 17 39 5.47996 $w=1.3e-08 $l=2.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1160 $X2=0.6210 $Y2=0.1395
r27 37 38 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1530 $X2=0.2045 $Y2=0.1530
r28 37 45 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1890 $Y=0.1530
+ $X2=0.1890 $Y2=0.1530
r29 35 38 16.2067 $w=1.3e-08 $l=6.95e-08 $layer=M2 $thickness=3.6e-08 $X=0.2740
+ $Y=0.1530 $X2=0.2045 $Y2=0.1530
r30 33 34 15.2739 $w=1.3e-08 $l=6.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1530 $X2=0.6865 $Y2=0.1530
r31 33 39 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.6210 $Y=0.1530 $X2=0.6210
+ $Y2=0.1395
r32 32 33 34.1623 $w=1.3e-08 $l=1.465e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.4745 $Y=0.1530 $X2=0.6210 $Y2=0.1530
r33 32 35 46.7545 $w=1.3e-08 $l=2.005e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.4745 $Y=0.1530 $X2=0.2740 $Y2=0.1530
r34 22 31 18.3054 $w=1.3e-08 $l=7.85e-08 $layer=M2 $thickness=3.6e-08 $X=0.8125
+ $Y=0.1530 $X2=0.8910 $Y2=0.1530
r35 22 34 29.3819 $w=1.3e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.8125
+ $Y=0.1530 $X2=0.6865 $Y2=0.1530
r36 29 31 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.8910 $Y=0.1440
+ $X2=0.8910 $Y2=0.1530
r37 18 29 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1135 $X2=0.8910 $Y2=0.1440
r38 12 2 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.8910
+ $Y=0.1350 $X2=0.8910 $Y2=0.1350
r39 2 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8910 $Y=0.1350
+ $X2=0.8910 $Y2=0.1440
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%SH VSS 11 12 13 75 78 80 83 15 16 22 24 14 6 19
+ 17 18 5 21 2 26 23 1 20 25
c1 1 VSS 0.000629939f
c2 2 VSS 0.00773759f
c3 5 VSS 0.0049912f
c4 6 VSS 0.00514847f
c5 11 VSS 0.0377083f
c6 12 VSS 0.0807875f
c7 13 VSS 0.0809773f
c8 14 VSS 0.00514527f
c9 15 VSS 0.00531115f
c10 16 VSS 0.00800877f
c11 17 VSS 0.000583789f
c12 18 VSS 0.00159113f
c13 19 VSS 0.0012234f
c14 20 VSS 0.000162985f
c15 21 VSS 0.00493712f
c16 22 VSS 0.00673915f
c17 23 VSS 0.00221217f
c18 24 VSS 0.000166949f
c19 25 VSS 0.000430893f
c20 26 VSS 0.0158968f
r1 83 82 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8810 $Y=0.0405 $X2=0.8785 $Y2=0.0405
r2 5 82 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8660 $Y=0.0405 $X2=0.8785 $Y2=0.0405
r3 79 5 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8540 $Y=0.0405 $X2=0.8660 $Y2=0.0405
r4 14 79 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.0405 $X2=0.8540 $Y2=0.0405
r5 80 14 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.0405 $X2=0.8495 $Y2=0.0405
r6 78 77 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9350 $Y=0.2295 $X2=0.9325 $Y2=0.2295
r7 76 77 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9280 $Y=0.2295 $X2=0.9325 $Y2=0.2295
r8 6 76 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9160 $Y=0.2295 $X2=0.9280 $Y2=0.2295
r9 15 6 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9035 $Y=0.2295 $X2=0.9160 $Y2=0.2295
r10 75 15 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9010 $Y=0.2295 $X2=0.9035 $Y2=0.2295
r11 13 68 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=1.3230
+ $Y=0.1350 $X2=1.3230 $Y2=0.1360
r12 12 60 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=1.2690 $Y=0.1350 $X2=1.2690 $Y2=0.1360
r13 5 58 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.0405
+ $X2=0.8640 $Y2=0.0360
r14 6 53 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.9180 $Y=0.2295
+ $X2=0.9180 $Y2=0.2340
r15 66 68 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.3105 $Y=0.1360 $X2=1.3230 $Y2=0.1360
r16 65 66 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.2960 $Y=0.1360 $X2=1.3105 $Y2=0.1360
r17 63 65 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.2815 $Y=0.1360 $X2=1.2960 $Y2=0.1360
r18 61 63 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=1.2785 $Y=0.1360 $X2=1.2815 $Y2=0.1360
r19 60 61 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=1.2690
+ $Y=0.1360 $X2=1.2785 $Y2=0.1360
r20 2 60 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=1.2595
+ $Y=0.1360 $X2=1.2690 $Y2=0.1360
r21 58 59 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.0360 $X2=0.8775 $Y2=0.0360
r22 56 59 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.0360 $X2=0.8775 $Y2=0.0360
r23 55 56 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.9020
+ $Y=0.0360 $X2=0.8910 $Y2=0.0360
r24 16 23 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.9200
+ $Y=0.0360 $X2=0.9450 $Y2=0.0360
r25 16 55 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.9200
+ $Y=0.0360 $X2=0.9020 $Y2=0.0360
r26 53 54 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.2340 $X2=0.9315 $Y2=0.2340
r27 22 54 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.2340 $X2=0.9315 $Y2=0.2340
r28 50 60 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.2690 $Y=0.1445
+ $X2=1.2690 $Y2=0.1360
r29 21 50 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.2690
+ $Y=0.1085 $X2=1.2690 $Y2=0.1445
r30 23 44 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.0360 $X2=0.9450 $Y2=0.0630
r31 18 39 6.50021 $w=1.33448e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.1980 $X2=0.9450 $Y2=0.1690
r32 18 22 7.21452 $w=1.425e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.1980 $X2=0.9450 $Y2=0.2340
r33 48 50 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=1.2690 $Y=0.1530
+ $X2=1.2690 $Y2=0.1445
r34 47 48 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=1.2445
+ $Y=0.1530 $X2=1.2690 $Y2=0.1530
r35 46 47 9.91056 $w=1.3e-08 $l=4.25e-08 $layer=M2 $thickness=3.6e-08 $X=1.2020
+ $Y=0.1530 $X2=1.2445 $Y2=0.1530
r36 45 46 32.0636 $w=1.3e-08 $l=1.375e-07 $layer=M2 $thickness=3.6e-08
+ $X=1.0645 $Y=0.1530 $X2=1.2020 $Y2=0.1530
r37 26 45 27.8662 $w=1.3e-08 $l=1.195e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.9450 $Y=0.1530 $X2=1.0645 $Y2=0.1530
r38 26 40 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.9450 $Y=0.1530 $X2=0.9450
+ $Y2=0.1485
r39 43 44 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.0900 $X2=0.9450 $Y2=0.0630
r40 42 43 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1000 $X2=0.9450 $Y2=0.0900
r41 41 42 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1100 $X2=0.9450 $Y2=0.1000
r42 17 40 3.96423 $w=1.3e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1315 $X2=0.9450 $Y2=0.1485
r43 17 41 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1315 $X2=0.9450 $Y2=0.1100
r44 38 39 0.4592 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1645 $X2=0.9450 $Y2=0.1690
r45 24 38 0.714311 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1575 $X2=0.9450 $Y2=0.1645
r46 24 40 1.50855 $w=1.55e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1575 $X2=0.9450 $Y2=0.1485
r47 24 26 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.9450 $Y=0.1575 $X2=0.9450
+ $Y2=0.1530
r48 37 39 4.4015 $w=1.35e-08 $l=2.78927e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9720 $Y=0.1620 $X2=0.9450 $Y2=0.1690
r49 36 37 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9990
+ $Y=0.1620 $X2=0.9720 $Y2=0.1620
r50 19 25 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0260 $Y=0.1620 $X2=1.0530 $Y2=0.1620
r51 19 36 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.1620 $X2=0.9990 $Y2=0.1620
r52 25 34 0.915974 $w=2.10182e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0530 $Y=0.1620 $X2=1.0530 $Y2=0.1510
r53 33 34 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1400 $X2=1.0530 $Y2=0.1510
r54 20 33 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1250 $X2=1.0530 $Y2=0.1400
r55 1 30 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=1.0530
+ $Y=0.1400 $X2=1.0530 $Y2=0.1400
r56 1 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.0530 $Y=0.1400
+ $X2=1.0530 $Y2=0.1400
r57 11 30 0.314665 $w=2.27e-07 $l=5e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.0530 $Y=0.1350 $X2=1.0530 $Y2=0.1400
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%CLKN VSS 16 17 18 19 20 101 103 30 27 26 31 8 22
+ 21 33 9 1 35 25 23 2 28 34 10 5 29 3 32 24
c1 1 VSS 0.00150475f
c2 2 VSS 0.000252022f
c3 3 VSS 5.45542e-20
c4 4 VSS 1e-36
c5 5 VSS 0.000278849f
c6 8 VSS 0.00776309f
c7 9 VSS 0.0080002f
c8 10 VSS 0.00382925f
c9 16 VSS 0.0593151f
c10 17 VSS 0.00583263f
c11 18 VSS 0.0050807f
c12 19 VSS 0.00437437f
c13 20 VSS 0.00534271f
c14 21 VSS 0.00645277f
c15 22 VSS 0.00637189f
c16 23 VSS 0.00789362f
c17 24 VSS 0.00177755f
c18 25 VSS 0.0046317f
c19 26 VSS 0.00375884f
c20 27 VSS 0.00114498f
c21 28 VSS 0.0025213f
c22 29 VSS 0.00137889f
c23 30 VSS 0.00366164f
c24 31 VSS 0.00197191f
c25 32 VSS 0.00396323f
c26 33 VSS 0.00138106f
c27 34 VSS 0.000587872f
c28 35 VSS 0.0298631f
r1 103 102 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r2 22 102 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r3 101 100 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r4 21 100 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r5 9 98 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0550 $Y2=0.2340
r6 8 95 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0550 $Y2=0.0360
r7 97 98 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.2340 $X2=0.0550 $Y2=0.2340
r8 26 97 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0460 $Y2=0.2340
r9 26 32 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0180 $Y2=0.2340
r10 94 95 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.0360 $X2=0.0550 $Y2=0.0360
r11 25 94 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0460 $Y2=0.0360
r12 25 30 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0180 $Y2=0.0360
r13 32 92 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.2340 $X2=0.0180 $Y2=0.2160
r14 30 91 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.0360 $X2=0.0180 $Y2=0.0630
r15 1 83 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
r16 16 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r17 24 31 1.81469 $w=1.6125e-08 $l=1.35831e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.2025 $X2=0.0165 $Y2=0.1890
r18 24 92 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.2025 $X2=0.0180 $Y2=0.2160
r19 90 91 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0900 $X2=0.0180 $Y2=0.0630
r20 89 90 9.67737 $w=1.3e-08 $l=4.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1315 $X2=0.0180 $Y2=0.0900
r21 23 31 2.63085 $w=1.54194e-08 $l=1.7066e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1720 $X2=0.0165 $Y2=0.1890
r22 23 89 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1720 $X2=0.0180 $Y2=0.1315
r23 2 74 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1355
+ $X2=0.5670 $Y2=0.1350
r24 17 2 3.19489 $w=1.24e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1355
r25 33 69 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.1350 $Y=0.1980 $X2=0.1350
+ $Y2=0.1890
r26 83 84 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1540
r27 81 84 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1720 $X2=0.1350 $Y2=0.1540
r28 27 69 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.1350 $Y=0.1845 $X2=0.1350
+ $Y2=0.1890
r29 27 81 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1845 $X2=0.1350 $Y2=0.1720
r30 27 33 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1845 $X2=0.1350 $Y2=0.1980
r31 78 79 1.90199 $w=1.38333e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.0255 $Y=0.1890 $X2=0.0345 $Y2=0.1890
r32 31 78 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0165
+ $Y=0.1890 $X2=0.0255 $Y2=0.1890
r33 34 71 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.1980 $X2=0.5670 $Y2=0.1845
r34 34 62 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.5670 $Y=0.1980 $X2=0.5670
+ $Y2=0.1890
r35 74 75 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1485
r36 72 75 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1620 $X2=0.5670 $Y2=0.1485
r37 28 71 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1755 $X2=0.5670 $Y2=0.1845
r38 28 72 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1755 $X2=0.5670 $Y2=0.1620
r39 69 70 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1890 $X2=0.1595 $Y2=0.1890
r40 68 69 11.8927 $w=1.3e-08 $l=5.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.0840
+ $Y=0.1890 $X2=0.1350 $Y2=0.1890
r41 67 68 11.8927 $w=1.3e-08 $l=5.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.0330
+ $Y=0.1890 $X2=0.0840 $Y2=0.1890
r42 67 79 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.0330 $Y=0.1890
+ $X2=0.0345 $Y2=0.1890
r43 63 64 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.6480
+ $Y=0.1890 $X2=0.7290 $Y2=0.1890
r44 62 63 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1890 $X2=0.6480 $Y2=0.1890
r45 62 71 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.5670 $Y=0.1890 $X2=0.5670
+ $Y2=0.1845
r46 35 62 46.7546 $w=1.3e-08 $l=2.005e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.3665 $Y=0.1890 $X2=0.5670 $Y2=0.1890
r47 35 70 48.2703 $w=1.3e-08 $l=2.07e-07 $layer=M2 $thickness=3.6e-08 $X=0.3665
+ $Y=0.1890 $X2=0.1595 $Y2=0.1890
r48 5 59 2.78395 $w=2.4e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.9450
+ $Y=0.1780 $X2=0.9450 $Y2=0.1780
r49 20 5 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.9450 $Y=0.1350 $X2=0.9450 $Y2=0.1780
r50 3 52 2.78395 $w=2.4e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.6750
+ $Y=0.1780 $X2=0.6750 $Y2=0.1780
r51 18 3 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.6750 $Y=0.1350 $X2=0.6750 $Y2=0.1780
r52 60 64 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.7290 $Y=0.1845
+ $X2=0.7290 $Y2=0.1890
r53 29 60 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1680 $X2=0.7290 $Y2=0.1845
r54 58 59 6.83711 $w=2.22e-08 $l=1.5e-09 $layer=LISD $thickness=2.7e-08
+ $X=0.9435 $Y=0.1780 $X2=0.9450 $Y2=0.1780
r55 57 58 12.9145 $w=2.22e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9180 $Y=0.1780 $X2=0.9435 $Y2=0.1780
r56 56 57 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9045 $Y=0.1780 $X2=0.9180 $Y2=0.1780
r57 55 56 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8910 $Y=0.1780 $X2=0.9045 $Y2=0.1780
r58 54 55 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8775 $Y=0.1780 $X2=0.8910 $Y2=0.1780
r59 53 54 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8640 $Y=0.1780 $X2=0.8775 $Y2=0.1780
r60 51 52 12.9145 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6885 $Y=0.1780 $X2=0.6750 $Y2=0.1780
r61 50 51 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7155 $Y=0.1780 $X2=0.6885 $Y2=0.1780
r62 48 49 6.07743 $w=2.22e-08 $l=1.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7290 $Y=0.1780 $X2=0.7410 $Y2=0.1780
r63 48 60 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7290 $Y=0.1780
+ $X2=0.7290 $Y2=0.1845
r64 47 48 5.31775 $w=2.22e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7185 $Y=0.1780 $X2=0.7290 $Y2=0.1780
r65 47 50 1.51936 $w=2.22e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.7185
+ $Y=0.1780 $X2=0.7155 $Y2=0.1780
r66 46 49 4.55807 $w=2.22e-08 $l=9e-09 $layer=LISD $thickness=2.7e-08 $X=0.7500
+ $Y=0.1780 $X2=0.7410 $Y2=0.1780
r67 45 46 6.07743 $w=2.22e-08 $l=1.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7620 $Y=0.1780 $X2=0.7500 $Y2=0.1780
r68 44 45 4.05162 $w=2.22e-08 $l=8e-09 $layer=LISD $thickness=2.7e-08 $X=0.7700
+ $Y=0.1780 $X2=0.7620 $Y2=0.1780
r69 43 44 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7835 $Y=0.1780 $X2=0.7700 $Y2=0.1780
r70 42 43 6.58388 $w=2.22e-08 $l=1.3e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7965 $Y=0.1780 $X2=0.7835 $Y2=0.1780
r71 41 42 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8100 $Y=0.1780 $X2=0.7965 $Y2=0.1780
r72 10 41 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8370 $Y=0.1780 $X2=0.8100 $Y2=0.1780
r73 10 53 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8370 $Y=0.1780 $X2=0.8640 $Y2=0.1780
r74 4 40 2.78395 $w=2.4e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.8370
+ $Y=0.1780 $X2=0.8370 $Y2=0.1780
r75 4 10 10.3807 $w=2.30357e-08 $l=0 $layer=LISD $thickness=3.675e-08 $X=0.8370
+ $Y=0.1780 $X2=0.8370 $Y2=0.1780
r76 19 40 0.314665 $w=2.27e-07 $l=4.3e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.8370 $Y=0.1350 $X2=0.8370 $Y2=0.1780
r77 9 22 1e-05
r78 8 21 1e-05
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%noxref_26 VSS 1
c1 1 VSS 0.00432565f
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%SI VSS 14 3 5 6 7 1 4
c1 1 VSS 0.00578422f
c2 3 VSS 0.00731476f
c3 4 VSS 0.00310641f
c4 5 VSS 0.00300212f
c5 6 VSS 0.00356204f
c6 7 VSS 0.00369797f
r1 6 19 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1980 $X2=0.5130 $Y2=0.1765
r2 5 7 3.2503 $w=1.53684e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1540 $X2=0.5130 $Y2=0.1350
r3 5 19 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1540 $X2=0.5130 $Y2=0.1765
r4 7 16 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1350 $X2=0.4945 $Y2=0.1350
r5 15 16 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4845
+ $Y=0.1350 $X2=0.4945 $Y2=0.1350
r6 14 15 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4750
+ $Y=0.1350 $X2=0.4845 $Y2=0.1350
r7 14 4 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4750
+ $Y=0.1350 $X2=0.4635 $Y2=0.1350
r8 14 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4750 $Y=0.1350
+ $X2=0.4790 $Y2=0.1350
r9 11 12 4.43042 $w=1.53e-08 $l=7.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.4715
+ $Y=0.1350 $X2=0.4790 $Y2=0.1350
r10 9 11 1.86855 $w=1.78125e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.4675 $Y=0.1350 $X2=0.4715 $Y2=0.1350
r11 1 9 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.4575
+ $Y=0.1350 $X2=0.4675 $Y2=0.1350
r12 3 1 2.53453 $w=1.32811e-07 $l=1.5e-09 $layer=LIG $thickness=5.23243e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4575 $Y2=0.1350
r13 3 11 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4715 $Y2=0.1350
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%noxref_28 VSS 1
c1 1 VSS 0.00573776f
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%noxref_30 VSS 1
c1 1 VSS 0.0124611f
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%NET0167 VSS 14 27 7 9 1 11 12 10 8 2
c1 1 VSS 0.00639051f
c2 2 VSS 0.00558077f
c3 7 VSS 0.00468324f
c4 8 VSS 0.00321658f
c5 9 VSS 0.000875426f
c6 10 VSS 0.0175502f
c7 11 VSS 0.00131907f
c8 12 VSS 0.0020732f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0675 $X2=0.4840 $Y2=0.0675
r2 27 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4715 $Y2=0.0675
r3 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0675
+ $X2=0.4860 $Y2=0.0360
r4 23 24 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4475
+ $Y=0.0360 $X2=0.4860 $Y2=0.0360
r5 22 23 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4070
+ $Y=0.0360 $X2=0.4475 $Y2=0.0360
r6 21 22 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.3875
+ $Y=0.0360 $X2=0.4070 $Y2=0.0360
r7 20 21 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3605
+ $Y=0.0360 $X2=0.3875 $Y2=0.0360
r8 19 20 7.92845 $w=1.3e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3265
+ $Y=0.0360 $X2=0.3605 $Y2=0.0360
r9 10 12 1.03257 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3085 $Y=0.0360 $X2=0.2970 $Y2=0.0360
r10 10 19 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3085
+ $Y=0.0360 $X2=0.3265 $Y2=0.0360
r11 12 18 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.2970 $Y2=0.0540
r12 9 17 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0720 $X2=0.2970 $Y2=0.0900
r13 9 18 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0720 $X2=0.2970 $Y2=0.0540
r14 16 17 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2835 $Y=0.0900 $X2=0.2970 $Y2=0.0900
r15 11 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0900 $X2=0.2835 $Y2=0.0900
r16 11 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0900
+ $X2=0.2700 $Y2=0.0945
r17 1 15 23.8708 $w=2.02e-08 $l=4.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.2700 $Y=0.0540 $X2=0.2700 $Y2=0.0945
r18 14 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r19 7 13 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r20 1 7 1e-05
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%PD1 VSS 12 13 29 8 2 9 7 1
c1 1 VSS 0.00351035f
c2 2 VSS 0.00381061f
c3 7 VSS 0.00294238f
c4 8 VSS 0.00227488f
c5 9 VSS 0.00244063f
r1 29 28 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.0675 $X2=0.6085 $Y2=0.0675
r2 27 28 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6040 $Y=0.0675 $X2=0.6085 $Y2=0.0675
r3 8 27 0.123457 $w=8.1e-08 $l=1e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.0675 $X2=0.6040 $Y2=0.0675
r4 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0675
+ $X2=0.5900 $Y2=0.0720
r5 23 24 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.5805
+ $Y=0.0720 $X2=0.5900 $Y2=0.0720
r6 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0720 $X2=0.5805 $Y2=0.0720
r7 21 22 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.0720 $X2=0.5670 $Y2=0.0720
r8 20 21 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0720 $X2=0.5400 $Y2=0.0720
r9 19 20 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5020
+ $Y=0.0720 $X2=0.5130 $Y2=0.0720
r10 18 19 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4805
+ $Y=0.0720 $X2=0.5020 $Y2=0.0720
r11 17 18 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.4540
+ $Y=0.0720 $X2=0.4805 $Y2=0.0720
r12 16 17 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4440
+ $Y=0.0720 $X2=0.4540 $Y2=0.0720
r13 15 16 1.63233 $w=1.3e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.4370
+ $Y=0.0720 $X2=0.4440 $Y2=0.0720
r14 14 15 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4280
+ $Y=0.0720 $X2=0.4370 $Y2=0.0720
r15 9 14 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4205
+ $Y=0.0720 $X2=0.4280 $Y2=0.0720
r16 1 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4280 $Y2=0.0720
r17 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r18 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r19 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0675 $X2=0.4320 $Y2=0.0675
r20 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4175 $Y2=0.0675
r21 2 8 1e-05
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%SE VSS 33 5 6 9 13 8 12 1 2 10 7 11
c1 1 VSS 0.00185327f
c2 2 VSS 0.0037858f
c3 5 VSS 0.0426606f
c4 6 VSS 0.0802896f
c5 7 VSS 0.00166985f
c6 8 VSS 0.000574275f
c7 9 VSS 0.0044862f
c8 10 VSS 0.00510911f
c9 11 VSS 0.00124536f
c10 12 VSS 0.00597839f
c11 13 VSS 0.0529809f
r1 1 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
r2 5 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r3 37 38 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2745
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r4 36 37 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2595
+ $Y=0.1350 $X2=0.2745 $Y2=0.1350
r5 35 36 0.699569 $w=1.3e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.1350 $X2=0.2595 $Y2=0.1350
r6 33 8 2.49951 $w=7.46154e-09 $l=1.95256e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.1340 $X2=0.2445 $Y2=0.1350
r7 8 35 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2445
+ $Y=0.1350 $X2=0.2565 $Y2=0.1350
r8 33 11 0.433689 $w=1.8e-08 $l=4.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.1340 $X2=0.2250 $Y2=0.1297
r9 11 31 3.53073 $w=1.4087e-08 $l=1.72e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.1297 $X2=0.2250 $Y2=0.1125
r10 10 27 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.2250 $Y=0.0360 $X2=0.2250
+ $Y2=0.0450
r11 30 31 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0900 $X2=0.2250 $Y2=0.1125
r12 29 30 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0675 $X2=0.2250 $Y2=0.0900
r13 7 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0495 $X2=0.2250 $Y2=0.0675
r14 7 27 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.2250 $Y=0.0495 $X2=0.2250
+ $Y2=0.0450
r15 7 10 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.0495 $X2=0.2250 $Y2=0.0360
r16 27 28 14.108 $w=1.3e-08 $l=6.05e-08 $layer=M2 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0450 $X2=0.2855 $Y2=0.0450
r17 25 28 109.716 $w=1.3e-08 $l=4.705e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.7560 $Y=0.0450 $X2=0.2855 $Y2=0.0450
r18 13 23 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=1.1905
+ $Y=0.0450 $X2=1.2150 $Y2=0.0450
r19 13 25 101.321 $w=1.3e-08 $l=4.345e-07 $layer=M2 $thickness=3.6e-08
+ $X=1.1905 $Y=0.0450 $X2=0.7560 $Y2=0.0450
r20 12 23 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=1.2150 $Y=0.0360 $X2=1.2150
+ $Y2=0.0450
r21 19 20 6.41272 $w=1.3e-08 $l=2.75e-08 $layer=M1 $thickness=3.6e-08 $X=1.2150
+ $Y=0.1085 $X2=1.2150 $Y2=0.1360
r22 18 19 8.51143 $w=1.3e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=1.2150
+ $Y=0.0720 $X2=1.2150 $Y2=0.1085
r23 9 18 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.2150
+ $Y=0.0495 $X2=1.2150 $Y2=0.0720
r24 9 12 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.2150 $Y=0.0495 $X2=1.2150 $Y2=0.0360
r25 9 23 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=1.2150 $Y=0.0495 $X2=1.2150
+ $Y2=0.0450
r26 17 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.2150 $Y=0.1380
+ $X2=1.2150 $Y2=0.1360
r27 6 2 1.49611 $w=1.91717e-07 $l=8e-09 $layer=LIG $thickness=5.46667e-08
+ $X=1.2150 $Y=0.1350 $X2=1.2150 $Y2=0.1270
r28 6 17 5.63117 $w=1.26721e-07 $l=3e-09 $layer=LIG $thickness=5.22105e-08
+ $X=1.2150 $Y=0.1350 $X2=1.2150 $Y2=0.1380
.ends

.subckt PM_SDFLx2_ASAP7_75t_R%SEN VSS 9 45 50 3 4 13 14 1 15 11 10 12 16
c1 1 VSS 0.00390895f
c2 3 VSS 0.0093204f
c3 4 VSS 0.00817242f
c4 9 VSS 0.081597f
c5 10 VSS 0.00503839f
c6 11 VSS 0.00534057f
c7 12 VSS 0.00167154f
c8 13 VSS 0.00333134f
c9 14 VSS 0.000818549f
c10 15 VSS 0.00580069f
c11 16 VSS 0.0131431f
r1 50 49 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.2050 $Y=0.2025 $X2=1.2025 $Y2=0.2025
r2 11 49 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.1900 $Y=0.2025 $X2=1.2025 $Y2=0.2025
r3 4 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.1880 $Y=0.2295
+ $X2=1.1880 $Y2=0.2340
r4 45 44 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.2050 $Y=0.0675 $X2=1.2025 $Y2=0.0675
r5 10 44 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.1900 $Y=0.0675 $X2=1.2025 $Y2=0.0675
r6 41 42 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.1745
+ $Y=0.2340 $X2=1.1880 $Y2=0.2340
r7 15 37 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1610 $Y=0.2340 $X2=1.1610 $Y2=0.2125
r8 15 41 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1610 $Y=0.2340 $X2=1.1745 $Y2=0.2340
r9 3 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.1725 $Y=0.0405
+ $X2=1.1610 $Y2=0.0515
r10 3 10 4.30736 $w=5.12e-08 $l=2.95e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.1725 $Y=0.0405 $X2=1.1725 $Y2=0.0700
r11 36 37 15.7403 $w=1.3e-08 $l=6.75e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.1450 $X2=1.1610 $Y2=0.2125
r12 35 36 14.9241 $w=1.3e-08 $l=6.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0810 $X2=1.1610 $Y2=0.1450
r13 34 35 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0650 $X2=1.1610 $Y2=0.0810
r14 33 34 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0515 $X2=1.1610 $Y2=0.0650
r15 32 33 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0425 $X2=1.1610 $Y2=0.0515
r16 13 32 1.28254 $w=1.3e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0370 $X2=1.1610 $Y2=0.0425
r17 30 35 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=1.1610 $Y=0.0810
+ $X2=1.1610 $Y2=0.0810
r18 29 30 27.2832 $w=1.3e-08 $l=1.17e-07 $layer=M2 $thickness=3.6e-08 $X=1.0440
+ $Y=0.0810 $X2=1.1610 $Y2=0.0810
r19 28 29 29.3819 $w=1.3e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.9180
+ $Y=0.0810 $X2=1.0440 $Y2=0.0810
r20 27 28 67.1587 $w=1.3e-08 $l=2.88e-07 $layer=M2 $thickness=3.6e-08 $X=0.6300
+ $Y=0.0810 $X2=0.9180 $Y2=0.0810
r21 26 27 65.0599 $w=1.3e-08 $l=2.79e-07 $layer=M2 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0810 $X2=0.6300 $Y2=0.0810
r22 16 26 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.3395
+ $Y=0.0810 $X2=0.3510 $Y2=0.0810
r23 14 22 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.0720 $X2=0.3510 $Y2=0.0855
r24 14 26 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.3510 $Y=0.0720 $X2=0.3510
+ $Y2=0.0810
r25 22 23 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0855 $X2=0.3510 $Y2=0.0945
r26 22 26 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.3510 $Y=0.0855 $X2=0.3510
+ $Y2=0.0810
r27 21 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1080 $X2=0.3510 $Y2=0.0945
r28 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1215 $X2=0.3510 $Y2=0.1080
r29 12 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1215
r30 9 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r31 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
r32 4 11 1e-05
.ends


*
.SUBCKT SDFLx2_ASAP7_75t_R VSS VDD CLK SE D SI QN
*
* VSS VSS
* VDD VDD
* CLK CLK
* SE SE
* D D
* SI SI
* QN QN
*
*

MM20 N_MM20_d N_MM20_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM23 N_MM23_d N_MM22_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM26 N_MM26_d N_MM31_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM29 N_MM29_d N_MM27_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM32 N_MM32_d N_MM30_g N_MM32_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM3_g N_MM5_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM10_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM6 N_MM6_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM12 N_MM12_d N_MM12_g N_MM12_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM17 N_MM17_d N_MM17_g N_MM17_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM16 N_MM16_d N_MM16_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM14 N_MM14_d N_MM14_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM0 N_MM0_d N_MM0_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24 N_MM24_d N_MM24_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@2 N_MM24@2_d N_MM24@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM21 N_MM21_d N_MM20_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM22 N_MM22_d N_MM22_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM31 N_MM31_d N_MM31_g N_MM31_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM27 N_MM27_d N_MM27_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM30 N_MM30_d N_MM30_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g N_MM3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM13 N_MM13_d N_MM17_g N_MM13_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM18 N_MM18_d N_MM18_g N_MM18_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM19 N_MM19_d N_MM16_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM15 N_MM15_d N_MM14_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM2 N_MM2_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25 N_MM25_d N_MM24_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@2 N_MM25@2_d N_MM24@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "SDFLx2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "SDFLx2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_SDFLx2_ASAP7_75t_R%NET0168 VSS N_MM29_d N_MM32_s N_NET0168_1
+ PM_SDFLx2_ASAP7_75t_R%NET0168
cc_1 N_NET0168_1 N_MM27_g 0.0173504f
cc_2 N_NET0168_1 N_MM30_g 0.0172405f
x_PM_SDFLx2_ASAP7_75t_R%noxref_34 VSS N_noxref_34_1
+ PM_SDFLx2_ASAP7_75t_R%noxref_34
cc_3 N_noxref_34_1 N_MM0_g 0.00135619f
cc_4 N_noxref_34_1 N_SEN_3 0.000120195f
cc_5 N_noxref_34_1 N_SEN_4 0.000413325f
cc_6 N_noxref_34_1 N_SEN_11 0.037307f
cc_7 N_noxref_34_1 N_noxref_31_1 0.000463912f
cc_8 N_noxref_34_1 N_noxref_32_1 0.00775191f
cc_9 N_noxref_34_1 N_noxref_33_1 0.00120915f
x_PM_SDFLx2_ASAP7_75t_R%noxref_33 VSS N_noxref_33_1
+ PM_SDFLx2_ASAP7_75t_R%noxref_33
cc_10 N_noxref_33_1 N_MM0_g 0.00130553f
cc_11 N_noxref_33_1 N_SEN_3 0.00192718f
cc_12 N_noxref_33_1 N_SEN_10 0.0374892f
cc_13 N_noxref_33_1 N_noxref_31_1 0.00746202f
cc_14 N_noxref_33_1 N_noxref_32_1 0.000448944f
x_PM_SDFLx2_ASAP7_75t_R%D VSS D N_MM30_g N_D_1 N_D_5 PM_SDFLx2_ASAP7_75t_R%D
cc_15 N_MM30_g N_SEN_16 0.000481843f
cc_16 N_MM30_g N_SEN_1 0.000865616f
cc_17 N_D_1 N_SEN_1 0.00120732f
cc_18 N_D_5 N_SEN_14 0.00159242f
cc_19 N_D N_SEN_12 0.0021517f
cc_20 N_MM30_g N_MM27_g 0.00504614f
x_PM_SDFLx2_ASAP7_75t_R%PD3 VSS N_MM9_s N_MM8_d N_PD3_1
+ PM_SDFLx2_ASAP7_75t_R%PD3
cc_21 N_PD3_1 N_MM9_g 0.00777478f
cc_22 N_PD3_1 N_MM11_g 0.0078334f
x_PM_SDFLx2_ASAP7_75t_R%PD4 VSS N_MM18_s N_MM19_d N_PD4_1
+ PM_SDFLx2_ASAP7_75t_R%PD4
cc_23 N_PD4_1 N_MM18_g 0.00783215f
cc_24 N_PD4_1 N_MM16_g 0.00773625f
x_PM_SDFLx2_ASAP7_75t_R%NET0144 VSS N_MM31_s N_MM27_d N_MM30_d N_MM3_s
+ N_NET0144_9 N_NET0144_7 N_NET0144_1 N_NET0144_2 N_NET0144_8
+ PM_SDFLx2_ASAP7_75t_R%NET0144
cc_25 N_NET0144_9 N_CLKN_35 0.00296035f
cc_26 N_NET0144_7 N_SE_1 0.000976128f
cc_27 N_NET0144_9 N_SE_8 0.000729057f
cc_28 N_NET0144_1 N_MM31_g 0.00083414f
cc_29 N_NET0144_7 N_MM31_g 0.0328594f
cc_30 N_NET0144_7 N_SEN_1 0.000919032f
cc_31 N_NET0144_1 N_MM27_g 0.000850858f
cc_32 N_NET0144_9 N_SEN_12 0.00208069f
cc_33 N_NET0144_7 N_MM27_g 0.0329446f
cc_34 N_NET0144_2 N_MM30_g 0.000864139f
cc_35 N_NET0144_9 N_D 0.00224335f
cc_36 N_NET0144_8 N_MM30_g 0.0339625f
cc_37 N_NET0144_9 N_SI_4 0.00061549f
cc_38 N_NET0144_8 N_SI_1 0.000776145f
cc_39 N_NET0144_2 N_MM3_g 0.000815023f
cc_40 N_NET0144_8 N_MM3_g 0.0335001f
cc_41 N_NET0144_2 N_PU1_11 0.000546842f
cc_42 N_NET0144_7 N_PU1_8 0.00110342f
cc_43 N_NET0144_8 N_PU1_9 0.000553893f
cc_44 N_NET0144_1 N_PU1_11 0.000596543f
cc_45 N_NET0144_8 N_PU1_2 0.00129778f
cc_46 N_NET0144_2 N_PU1_2 0.00160893f
cc_47 N_NET0144_1 N_PU1_1 0.00302502f
cc_48 N_NET0144_9 N_PU1_11 0.0128284f
x_PM_SDFLx2_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_SDFLx2_ASAP7_75t_R%noxref_25
cc_49 N_noxref_25_1 N_MM20_g 0.00368232f
cc_50 N_noxref_25_1 N_CLKN_9 0.00053883f
cc_51 N_noxref_25_1 N_CLKN_8 4.38889e-20
cc_52 N_noxref_25_1 N_CLKN_32 5.43516e-20
cc_53 N_noxref_25_1 N_CLKN_24 7.69541e-20
cc_54 N_noxref_25_1 N_CLKN_31 9.32278e-20
cc_55 N_noxref_25_1 N_CLKN_23 0.000273916f
cc_56 N_noxref_25_1 N_CLKN_22 0.0275171f
cc_57 N_noxref_25_1 N_noxref_24_1 0.00204652f
x_PM_SDFLx2_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_SDFLx2_ASAP7_75t_R%noxref_24
cc_58 N_noxref_24_1 N_MM20_g 0.00368531f
cc_59 N_noxref_24_1 N_CLKN_31 3.2883e-20
cc_60 N_noxref_24_1 N_CLKN_8 0.000549624f
cc_61 N_noxref_24_1 N_CLKN_9 4.41927e-20
cc_62 N_noxref_24_1 N_CLKN_30 5.49094e-20
cc_63 N_noxref_24_1 N_CLKN_23 0.000386626f
cc_64 N_noxref_24_1 N_CLKN_21 0.0275607f
x_PM_SDFLx2_ASAP7_75t_R%PU1 VSS N_MM31_d N_MM3_d N_MM1_s N_PU1_10 N_PU1_2
+ N_PU1_11 N_PU1_8 N_PU1_1 N_PU1_9 PM_SDFLx2_ASAP7_75t_R%PU1
cc_65 N_PU1_10 N_CLKN_28 0.000382017f
cc_66 N_PU1_10 N_MM22_g 3.38266e-20
cc_67 N_PU1_10 N_CLKN_35 8.76711e-20
cc_68 N_PU1_10 N_CLKN_2 0.00101407f
cc_69 N_PU1_10 N_CLKN_34 0.000340792f
cc_70 N_PU1_2 N_MM1_g 0.00159178f
cc_71 N_PU1_11 N_CLKN_35 0.00340042f
cc_72 N_PU1_10 N_MM1_g 0.0339334f
cc_73 N_PU1_8 N_SE_8 0.000751981f
cc_74 N_PU1_8 N_SE_1 0.00100483f
cc_75 N_PU1_1 N_MM31_g 0.0013164f
cc_76 N_PU1_8 N_MM31_g 0.0341581f
cc_77 N_PU1_2 N_SI_5 0.000639681f
cc_78 N_PU1_9 N_SI_1 0.00143758f
cc_79 N_PU1_2 N_SI_6 0.00293904f
cc_80 N_PU1_11 N_SI_6 0.00314957f
cc_81 N_PU1_9 N_MM3_g 0.0350648f
cc_82 N_PU1_2 N_MH_3 0.00119002f
cc_83 N_PU1_2 N_MH_12 0.00291929f
x_PM_SDFLx2_ASAP7_75t_R%CLK VSS CLK N_MM20_g N_CLK_4 N_CLK_6 N_CLK_1 N_CLK_5
+ PM_SDFLx2_ASAP7_75t_R%CLK
x_PM_SDFLx2_ASAP7_75t_R%noxref_29 VSS N_noxref_29_1
+ PM_SDFLx2_ASAP7_75t_R%noxref_29
cc_84 N_noxref_29_1 N_MM31_g 0.00147391f
cc_85 N_noxref_29_1 N_CLKB_14 0.000676709f
cc_86 N_noxref_29_1 N_PU1_8 0.0360715f
cc_87 N_noxref_29_1 N_noxref_26_1 0.000466528f
cc_88 N_noxref_29_1 N_noxref_27_1 0.00771768f
cc_89 N_noxref_29_1 N_noxref_28_1 0.00123961f
x_PM_SDFLx2_ASAP7_75t_R%noxref_27 VSS N_noxref_27_1
+ PM_SDFLx2_ASAP7_75t_R%noxref_27
cc_90 N_noxref_27_1 N_CLKN_1 0.000129336f
cc_91 N_noxref_27_1 N_MM22_g 0.0034281f
cc_92 N_noxref_27_1 N_CLKB_6 0.000367361f
cc_93 N_noxref_27_1 N_CLKB_14 0.0271354f
cc_94 N_noxref_27_1 N_PU1_8 0.000589552f
cc_95 N_noxref_27_1 N_noxref_26_1 0.00148611f
x_PM_SDFLx2_ASAP7_75t_R%PD2 VSS N_MM10_s N_MM11_d N_PD2_4 N_PD2_5 N_PD2_1
+ PM_SDFLx2_ASAP7_75t_R%PD2
cc_96 N_PD2_4 N_CLKN_29 8.52631e-20
cc_97 N_PD2_4 N_CLKN_10 0.000126152f
cc_98 N_PD2_4 N_CLKN_3 0.000277563f
cc_99 N_PD2_5 N_CLKN_10 0.00167248f
cc_100 N_PD2_1 N_MM9_g 0.00209547f
cc_101 N_PD2_5 N_MM9_g 0.00734641f
cc_102 N_PD2_4 N_MM9_g 0.0237437f
cc_103 N_PD2_4 N_MM10_g 0.0150084f
cc_104 N_PD2_5 N_MM11_g 0.0148536f
cc_105 N_PD2_4 N_MH_14 0.000321594f
cc_106 N_PD2_4 N_MH_3 0.000612724f
cc_107 N_PD2_1 N_MH_14 0.00348294f
x_PM_SDFLx2_ASAP7_75t_R%noxref_35 VSS N_noxref_35_1
+ PM_SDFLx2_ASAP7_75t_R%noxref_35
cc_108 N_noxref_35_1 N_MM24@2_g 0.00148415f
cc_109 N_noxref_35_1 N_QN_7 0.000831772f
x_PM_SDFLx2_ASAP7_75t_R%noxref_32 VSS N_noxref_32_1
+ PM_SDFLx2_ASAP7_75t_R%noxref_32
cc_110 N_noxref_32_1 N_SEN_4 0.000150197f
cc_111 N_noxref_32_1 N_SEN_11 0.000893227f
cc_112 N_noxref_32_1 N_SS_11 0.0169645f
cc_113 N_noxref_32_1 N_MM14_g 0.0058046f
cc_114 N_noxref_32_1 N_noxref_31_1 0.00152625f
x_PM_SDFLx2_ASAP7_75t_R%noxref_31 VSS N_noxref_31_1
+ PM_SDFLx2_ASAP7_75t_R%noxref_31
cc_115 N_noxref_31_1 N_SEN_3 0.00180862f
cc_116 N_noxref_31_1 N_SS_10 0.0168945f
cc_117 N_noxref_31_1 N_MM14_g 0.00571276f
x_PM_SDFLx2_ASAP7_75t_R%SS VSS N_MM16_g N_MM14_d N_MM15_d N_SS_13 N_SS_15
+ N_SS_14 N_SS_17 N_SS_16 N_SS_12 N_SS_3 N_SS_4 N_SS_1 N_SS_10 N_SS_11
+ PM_SDFLx2_ASAP7_75t_R%SS
cc_118 N_MM16_g N_CLKN_10 0.000678009f
cc_119 N_MM16_g N_CLKN_5 0.000426619f
cc_120 N_MM16_g N_MM18_g 0.0133631f
cc_121 N_SS_13 N_SE_13 0.000905372f
cc_122 N_SS_15 N_SE_13 0.00323118f
cc_123 N_SS_14 N_SEN_3 0.00158892f
cc_124 N_SS_14 N_SEN_11 0.000118716f
cc_125 N_SS_14 N_SEN_15 0.000121753f
cc_126 N_SS_14 N_SEN_4 0.000255586f
cc_127 N_SS_13 N_SEN_16 0.000361395f
cc_128 N_SS_17 N_SEN_13 0.000429155f
cc_129 N_SS_16 N_SEN_15 0.000775661f
cc_130 N_SS_12 N_SEN_16 0.00262129f
cc_131 N_SS_14 N_SEN_13 0.00860387f
x_PM_SDFLx2_ASAP7_75t_R%noxref_36 VSS N_noxref_36_1
+ PM_SDFLx2_ASAP7_75t_R%noxref_36
cc_132 N_noxref_36_1 N_MM24@2_g 0.0014985f
cc_133 N_noxref_36_1 N_QN_8 0.000833507f
cc_134 N_noxref_36_1 N_noxref_35_1 0.00177631f
x_PM_SDFLx2_ASAP7_75t_R%PD5 VSS N_MM17_s N_MM16_d N_PD5_1 N_PD5_5 N_PD5_4
+ PM_SDFLx2_ASAP7_75t_R%PD5
cc_135 N_PD5_1 N_MM18_g 0.000757642f
cc_136 N_PD5_5 N_MM18_g 0.00693367f
cc_137 N_PD5_4 N_MM18_g 0.0239653f
cc_138 N_PD5_4 N_MM17_g 0.0152557f
cc_139 N_PD5_1 N_MM16_g 0.000892071f
cc_140 N_PD5_5 N_MM16_g 0.0155951f
cc_141 N_PD5_1 N_SH_14 0.000514906f
cc_142 N_PD5_1 N_SH_16 0.000490473f
cc_143 N_PD5_1 N_SH_17 0.000570926f
cc_144 N_PD5_4 N_SH_5 0.000658108f
cc_145 N_PD5_1 N_SH_23 0.0023807f
x_PM_SDFLx2_ASAP7_75t_R%QN VSS QN N_MM24_d N_MM24@2_d N_MM25_d N_MM25@2_d
+ N_QN_9 N_QN_7 N_QN_8 N_QN_10 N_QN_11 N_QN_1 N_QN_2 PM_SDFLx2_ASAP7_75t_R%QN
cc_146 N_QN_9 N_MM0_g 6.51622e-20
cc_147 N_QN_9 N_SE_9 0.000528237f
cc_148 N_QN_9 N_SE_13 0.000257635f
cc_149 N_QN_9 N_SE_12 0.00161575f
cc_150 N_QN_7 N_SH_21 0.000913751f
cc_151 N_QN_7 N_SH_2 0.000438658f
cc_152 N_QN_7 N_SH_26 0.000626074f
cc_153 N_QN_8 N_MM24_g 0.0308322f
cc_154 N_QN_10 N_SH_21 0.000951545f
cc_155 N_QN_11 N_SH_2 0.00118169f
cc_156 N_QN_1 N_MM24_g 0.00202951f
cc_157 N_QN_2 N_MM24_g 0.00241479f
cc_158 N_QN_2 N_SH_21 0.00259362f
cc_159 N_QN_8 N_SH_2 0.00471127f
cc_160 N_QN_7 N_MM24@2_g 0.0371529f
cc_161 N_QN_7 N_MM24_g 0.0682654f
x_PM_SDFLx2_ASAP7_75t_R%MH VSS N_MM7_g N_MM4_d N_MM9_d N_MM1_d N_MM10_d N_MH_10
+ N_MH_3 N_MH_21 N_MH_17 N_MH_1 N_MH_4 N_MH_12 N_MH_14 N_MH_18 N_MH_20 N_MH_16
+ N_MH_19 N_MH_15 PM_SDFLx2_ASAP7_75t_R%MH
cc_162 N_MH_10 N_CLKN_28 0.000122558f
cc_163 N_MH_10 N_CLKN_29 0.000340782f
cc_164 N_MH_10 N_MM1_g 0.000428002f
cc_165 N_MH_10 N_CLKN_2 0.000202873f
cc_166 N_MH_3 N_CLKN_28 0.000340115f
cc_167 N_MH_3 N_CLKN_34 0.000359138f
cc_168 N_MH_21 N_CLKN_29 0.000403742f
cc_169 N_MH_17 N_CLKN_29 0.00607883f
cc_170 N_MH_17 N_CLKN_3 0.000497072f
cc_171 N_MH_1 N_CLKN_10 0.00208388f
cc_172 N_MH_4 N_MM9_g 0.000633168f
cc_173 N_MH_12 N_CLKN_2 0.000667181f
cc_174 N_MH_17 N_CLKN_10 0.000773293f
cc_175 N_MH_14 N_CLKN_35 0.00141014f
cc_176 N_MH_18 N_CLKN_29 0.00149878f
cc_177 N_MH_3 N_MM1_g 0.00156222f
cc_178 N_MH_14 N_CLKN_34 0.00377168f
cc_179 N_MM7_g N_CLKN_10 0.00508184f
cc_180 N_MH_12 N_MM1_g 0.0329603f
cc_181 N_MM7_g N_MM12_g 0.0127275f
cc_182 N_MH_10 N_MM9_g 0.0361384f
cc_183 N_MH_10 N_CLKB_17 0.000251818f
cc_184 N_MH_10 N_CLKB_2 0.000109687f
cc_185 N_MH_10 N_MM17_g 0.000136903f
cc_186 N_MH_10 N_CLKB_21 0.000293692f
cc_187 N_MH_20 N_CLKB_21 0.00031856f
cc_188 N_MH_14 N_CLKB_21 0.000448847f
cc_189 N_MH_12 N_MM10_g 0.0163568f
cc_190 N_MH_16 N_CLKB_17 0.000526718f
cc_191 N_MH_3 N_CLKB_1 0.000604587f
cc_192 N_MH_4 N_CLKB_17 0.00080755f
cc_193 N_MH_4 N_MM10_g 0.00111037f
cc_194 N_MH_3 N_MM10_g 0.00122376f
cc_195 N_MH_10 N_CLKB_1 0.00160723f
cc_196 N_MH_17 N_CLKB_21 0.00205878f
cc_197 N_MH_18 N_CLKB_22 0.00250298f
cc_198 N_MH_10 N_MM10_g 0.0526632f
cc_199 N_MH_19 N_MS_18 0.000267048f
cc_200 N_MH_4 N_MS_1 0.00036012f
cc_201 N_MH_18 N_MS_19 0.000373635f
cc_202 N_MH_18 N_MS_1 0.000662301f
cc_203 N_MM7_g N_MS_3 0.000936962f
cc_204 N_MH_18 N_MS_17 0.000996507f
cc_205 N_MH_1 N_MS_14 0.00100248f
cc_206 N_MH_1 N_MS_1 0.0013014f
cc_207 N_MM7_g N_MS_12 0.00632007f
cc_208 N_MM7_g N_MS_1 0.00241085f
cc_209 N_MM7_g N_MS_11 0.00638981f
cc_210 N_MH_18 N_MS_14 0.00458906f
cc_211 N_MH_16 N_MS_18 0.00497056f
cc_212 N_MM7_g N_MM11_g 0.0293383f
x_PM_SDFLx2_ASAP7_75t_R%MS VSS N_MM11_g N_MM6_d N_MM12_d N_MM7_d N_MM13_d
+ N_MS_3 N_MS_15 N_MS_13 N_MS_12 N_MS_1 N_MS_17 N_MS_11 N_MS_4 N_MS_18 N_MS_19
+ N_MS_14 N_MS_16 PM_SDFLx2_ASAP7_75t_R%MS
cc_213 N_MS_3 N_CLKN_29 0.00014273f
cc_214 N_MS_3 N_CLKN_10 0.000652432f
cc_215 N_MS_3 N_CLKN_3 9.25654e-20
cc_216 N_MS_3 N_CLKN_35 0.000141518f
cc_217 N_MS_15 N_CLKN_29 0.000281055f
cc_218 N_MS_13 N_MM12_g 0.00786932f
cc_219 N_MS_15 N_CLKN_10 0.000361999f
cc_220 N_MS_12 N_MM12_g 0.00781547f
cc_221 N_MS_1 N_MM9_g 0.000704144f
cc_222 N_MS_17 N_CLKN_10 0.00154171f
cc_223 N_MS_11 N_MM12_g 0.006509f
cc_224 N_MS_4 N_MM12_g 0.00257216f
cc_225 N_MS_4 N_CLKN_10 0.00639182f
cc_226 N_MM11_g N_MM9_g 0.0141679f
cc_227 N_MS_3 N_MM12_g 0.0259814f
cc_228 N_MS_18 N_SEN_16 0.000922109f
cc_229 N_MS_19 N_SEN_16 0.00303756f
cc_230 N_MS_13 N_MM10_g 0.000137844f
cc_231 N_MS_13 N_CLKB_22 0.000349468f
cc_232 N_MS_13 N_CLKB_18 0.000180975f
cc_233 N_MS_13 N_CLKB_2 0.000222252f
cc_234 N_MS_17 N_CLKB_18 0.0045503f
cc_235 N_MS_17 N_CLKB_2 0.000289706f
cc_236 N_MS_19 N_CLKB_18 0.000418989f
cc_237 N_MS_18 N_CLKB_22 0.00167689f
cc_238 N_MS_13 N_MM17_g 0.0155691f
x_PM_SDFLx2_ASAP7_75t_R%CLKB VSS N_MM10_g N_MM17_g N_MM23_d N_MM22_d N_CLKB_13
+ N_CLKB_22 N_CLKB_16 N_CLKB_5 N_CLKB_19 N_CLKB_15 N_CLKB_6 N_CLKB_20 N_CLKB_14
+ N_CLKB_17 N_CLKB_18 N_CLKB_2 N_CLKB_1 N_CLKB_21 PM_SDFLx2_ASAP7_75t_R%CLKB
cc_239 N_CLKB_13 N_CLK_5 7.99986e-20
cc_240 N_CLKB_22 N_CLK_5 0.00012072f
cc_241 N_CLKB_16 N_CLK_5 0.000545769f
cc_242 N_CLKB_5 N_CLK_5 0.000386667f
cc_243 N_CLKB_19 N_CLK_5 0.00220898f
cc_244 N_CLKB_22 N_CLKN_10 2.85014e-20
cc_245 N_CLKB_22 N_CLKN_8 3.26977e-20
cc_246 N_CLKB_22 N_CLKN_25 3.59144e-20
cc_247 N_CLKB_22 N_MM22_g 4.9972e-20
cc_248 N_CLKB_5 N_CLKN_23 6.7653e-20
cc_249 N_CLKB_15 N_CLKN_26 0.00010366f
cc_250 N_CLKB_19 N_CLKN_27 0.000123067f
cc_251 N_CLKB_6 N_CLKN_33 0.000176973f
cc_252 N_MM17_g N_CLKN_5 0.000208159f
cc_253 N_CLKB_20 N_CLKN_33 0.000230779f
cc_254 N_CLKB_22 N_CLKN_29 0.000676953f
cc_255 N_CLKB_22 N_CLKN_28 0.000327609f
cc_256 N_CLKB_15 N_CLKN_27 0.000370527f
cc_257 N_CLKB_13 N_MM22_g 0.0386446f
cc_258 N_CLKB_14 N_MM22_g 0.0111649f
cc_259 N_CLKB_17 N_CLKN_35 0.000478614f
cc_260 N_CLKB_18 N_CLKN_10 0.000531969f
cc_261 N_CLKB_16 N_CLKN_1 0.000556157f
cc_262 N_MM10_g N_CLKN_3 0.000560153f
cc_263 N_CLKB_5 N_MM22_g 0.000594332f
cc_264 N_CLKB_16 N_CLKN_35 0.000617175f
cc_265 N_CLKB_2 N_CLKN_10 0.0027913f
cc_266 N_CLKB_14 N_CLKN_1 0.000776391f
cc_267 N_CLKB_6 N_MM22_g 0.000849536f
cc_268 N_CLKB_1 N_CLKN_2 0.00222254f
cc_269 N_CLKB_21 N_CLKN_34 0.00165668f
cc_270 N_CLKB_17 N_CLKN_28 0.00265567f
cc_271 N_CLKB_15 N_CLKN_33 0.00352324f
cc_272 N_MM10_g N_MM9_g 0.00370405f
cc_273 N_CLKB_16 N_CLKN_27 0.00487527f
cc_274 N_MM17_g N_CLKN_10 0.00493087f
cc_275 N_MM17_g N_MM18_g 0.00578278f
cc_276 N_MM10_g N_MM1_g 0.00704176f
cc_277 N_MM17_g N_MM12_g 0.0182753f
cc_278 N_CLKB_22 N_CLKN_35 0.0446295f
cc_279 N_CLKB_16 N_SE_1 5.26109e-20
cc_280 N_CLKB_5 N_SE_10 5.47477e-20
cc_281 N_CLKB_5 N_SE_7 0.000170428f
cc_282 N_CLKB_16 N_SE_7 0.00331576f
cc_283 N_CLKB_18 N_SE_13 0.000493925f
cc_284 N_CLKB_19 N_SE_10 0.00196725f
cc_285 N_CLKB_22 N_SE_13 0.00235535f
cc_286 N_CLKB_22 N_SE_8 0.00357527f
cc_287 N_CLKB_16 N_SE_11 0.00678176f
cc_288 N_CLKB_17 N_SEN_16 0.000503602f
cc_289 N_CLKB_22 N_SEN_12 0.00413661f
cc_290 N_CLKB_18 N_SEN_16 0.00281075f
cc_291 N_CLKB_22 N_SEN_16 0.00995479f
cc_292 N_CLKB_22 N_SI_4 0.00248603f
x_PM_SDFLx2_ASAP7_75t_R%SH VSS N_MM14_g N_MM24_g N_MM24@2_g N_MM13_s N_MM18_d
+ N_MM12_s N_MM17_d N_SH_15 N_SH_16 N_SH_22 N_SH_24 N_SH_14 N_SH_6 N_SH_19
+ N_SH_17 N_SH_18 N_SH_5 N_SH_21 N_SH_2 N_SH_26 N_SH_23 N_SH_1 N_SH_20 N_SH_25
+ PM_SDFLx2_ASAP7_75t_R%SH
cc_293 N_SH_15 N_CLKN_10 8.3963e-20
cc_294 N_SH_16 N_CLKN_35 9.21596e-20
cc_295 N_SH_22 N_CLKN_10 0.000196768f
cc_296 N_SH_24 N_CLKN_10 0.000203975f
cc_297 N_SH_14 N_MM12_g 0.00680288f
cc_298 N_SH_6 N_CLKN_10 0.000276295f
cc_299 N_SH_19 N_CLKN_10 0.000396208f
cc_300 N_SH_17 N_CLKN_10 0.000448364f
cc_301 N_SH_18 N_CLKN_10 0.000562805f
cc_302 N_SH_15 N_CLKN_5 0.000673075f
cc_303 N_SH_6 N_MM18_g 0.00100239f
cc_304 N_SH_5 N_CLKN_10 0.00282661f
cc_305 N_SH_5 N_MM12_g 0.00947937f
cc_306 N_SH_15 N_MM18_g 0.0160733f
cc_307 N_SH_21 N_SE_12 0.000231167f
cc_308 N_SH_17 N_SE_13 0.000315749f
cc_309 N_SH_2 N_SE_2 0.00163478f
cc_310 N_SH_16 N_SE_13 0.00102395f
cc_311 N_SH_26 N_SE_13 0.00209692f
cc_312 N_SH_23 N_SE_13 0.00268187f
cc_313 N_MM24_g N_MM0_g 0.00333059f
cc_314 N_SH_21 N_SE_9 0.00608386f
cc_315 N_MM24_g N_SEN_10 5.93708e-20
cc_316 N_SH_1 N_SEN_3 0.000208718f
cc_317 N_MM24_g N_SEN_4 0.000101615f
cc_318 N_SH_19 N_SEN_16 0.00010979f
cc_319 N_MM14_g N_SEN_3 0.000113039f
cc_320 N_SH_26 N_SEN_15 0.000117382f
cc_321 N_SH_26 N_SEN_13 0.00153856f
cc_322 N_SH_21 N_SEN_4 0.00019333f
cc_323 N_MM24_g N_SEN_3 0.000197376f
cc_324 N_SH_21 N_SEN_15 0.000261213f
cc_325 N_SH_20 N_SEN_16 0.000292155f
cc_326 N_SH_16 N_SEN_16 0.000373574f
cc_327 N_SH_26 N_SEN_16 0.00458679f
cc_328 N_SH_17 N_SEN_16 0.00609241f
cc_329 N_SH_6 N_MM17_g 0.000158318f
cc_330 N_SH_14 N_MM17_g 0.00676966f
cc_331 N_SH_15 N_MM17_g 0.00683991f
cc_332 N_SH_22 N_CLKB_18 0.000285306f
cc_333 N_SH_16 N_CLKB_18 0.000369687f
cc_334 N_SH_24 N_CLKB_18 0.000402567f
cc_335 N_SH_18 N_CLKB_18 0.000478333f
cc_336 N_SH_17 N_CLKB_2 0.000570191f
cc_337 N_SH_5 N_CLKB_2 0.000576027f
cc_338 N_SH_26 N_CLKB_22 0.000776466f
cc_339 N_SH_16 N_CLKB_22 0.0010628f
cc_340 N_SH_17 N_CLKB_18 0.00451947f
cc_341 N_SH_5 N_MM17_g 0.0183312f
cc_342 N_SH_18 N_MS_3 9.84546e-20
cc_343 N_SH_22 N_MS_3 0.000179155f
cc_344 N_SH_15 N_MS_3 0.000436412f
cc_345 N_SH_6 N_MS_3 0.000220896f
cc_346 N_SH_14 N_MS_3 0.000232021f
cc_347 N_SH_14 N_MS_11 0.000234022f
cc_348 N_SH_22 N_MS_4 0.000335655f
cc_349 N_SH_6 N_MS_4 0.000424812f
cc_350 N_SH_16 N_MS_16 0.00043823f
cc_351 N_SH_22 N_MS_17 0.000518125f
cc_352 N_SH_15 N_MS_4 0.00059315f
cc_353 N_SH_16 N_MS_19 0.00132439f
cc_354 N_SH_5 N_MS_3 0.00373419f
cc_355 N_SH_18 N_MM16_g 0.000104033f
cc_356 N_SH_20 N_SS_13 0.000310651f
cc_357 N_MM14_g N_SS_3 0.000322178f
cc_358 N_MM14_g N_SS_4 0.000425437f
cc_359 N_SH_23 N_SS_15 0.000580125f
cc_360 N_SH_25 N_SS_16 0.000623015f
cc_361 N_SH_25 N_SS_14 0.000697123f
cc_362 N_SH_17 N_SS_1 0.000810777f
cc_363 N_SH_1 N_SS_14 0.000950422f
cc_364 N_MM14_g N_SS_1 0.00111309f
cc_365 N_SH_1 N_MM16_g 0.00129928f
cc_366 N_SH_19 N_SS_12 0.00154842f
cc_367 N_SH_26 N_SS_14 0.00169853f
cc_368 N_MM14_g N_SS_10 0.00649523f
cc_369 N_MM14_g N_SS_11 0.00660041f
cc_370 N_SH_17 N_SS_12 0.00462671f
cc_371 N_SH_20 N_SS_14 0.00473501f
cc_372 N_MM14_g N_MM16_g 0.0300229f
x_PM_SDFLx2_ASAP7_75t_R%CLKN VSS N_MM22_g N_MM1_g N_MM9_g N_MM12_g N_MM18_g
+ N_MM20_d N_MM21_d N_CLKN_30 N_CLKN_27 N_CLKN_26 N_CLKN_31 N_CLKN_8 N_CLKN_22
+ N_CLKN_21 N_CLKN_33 N_CLKN_9 N_CLKN_1 N_CLKN_35 N_CLKN_25 N_CLKN_23 N_CLKN_2
+ N_CLKN_28 N_CLKN_34 N_CLKN_10 N_CLKN_5 N_CLKN_29 N_CLKN_3 N_CLKN_32 N_CLKN_24
+ PM_SDFLx2_ASAP7_75t_R%CLKN
cc_373 N_CLKN_30 N_MM20_g 5.92436e-20
cc_374 N_CLKN_27 N_MM20_g 7.17161e-20
cc_375 N_CLKN_26 N_MM20_g 8.98024e-20
cc_376 N_CLKN_31 N_MM20_g 9.82147e-20
cc_377 N_CLKN_8 N_MM20_g 0.00111234f
cc_378 N_CLKN_22 N_MM20_g 0.0112003f
cc_379 N_CLKN_21 N_MM20_g 0.0112112f
cc_380 N_CLKN_33 N_MM20_g 0.000355378f
cc_381 N_CLKN_31 N_CLK_4 0.000415112f
cc_382 N_CLKN_9 N_MM20_g 0.000630561f
cc_383 N_CLKN_1 N_CLK_6 0.00063244f
cc_384 N_CLKN_35 N_CLK_4 0.000647326f
cc_385 N_CLKN_25 N_CLK_6 0.000943393f
cc_386 N_CLKN_27 N_CLK_6 0.000948166f
cc_387 N_CLKN_1 N_CLK_1 0.00348994f
cc_388 N_CLKN_23 N_CLK_4 0.00164951f
cc_389 N_CLKN_25 N_CLK_5 0.00176865f
cc_390 N_CLKN_27 N_CLK_4 0.00477919f
cc_391 N_MM22_g N_MM20_g 0.0350676f
x_PM_SDFLx2_ASAP7_75t_R%noxref_26 VSS N_noxref_26_1
+ PM_SDFLx2_ASAP7_75t_R%noxref_26
cc_392 N_noxref_26_1 N_CLKN_1 0.000129154f
cc_393 N_noxref_26_1 N_MM22_g 0.00339694f
cc_394 N_noxref_26_1 N_CLKB_5 0.000434421f
cc_395 N_noxref_26_1 N_CLKB_13 0.0271823f
cc_396 N_noxref_26_1 N_NET0167_7 0.000552893f
x_PM_SDFLx2_ASAP7_75t_R%SI VSS SI N_MM3_g N_SI_5 N_SI_6 N_SI_7 N_SI_1 N_SI_4
+ PM_SDFLx2_ASAP7_75t_R%SI
cc_397 N_SI_5 N_CLKN_2 0.000464688f
cc_398 N_SI_5 N_MM1_g 7.57729e-20
cc_399 N_SI_5 N_CLKN_35 0.00103853f
cc_400 N_SI_6 N_CLKN_35 0.000321601f
cc_401 N_SI_7 N_CLKN_28 0.000820405f
cc_402 N_SI_6 N_CLKN_34 0.000920438f
cc_403 N_SI_5 N_CLKN_28 0.00259564f
cc_404 N_SI_1 N_MM30_g 0.000900113f
cc_405 N_SI_4 N_D_5 0.00100819f
cc_406 N_MM3_g N_MM30_g 0.00404453f
x_PM_SDFLx2_ASAP7_75t_R%noxref_28 VSS N_noxref_28_1
+ PM_SDFLx2_ASAP7_75t_R%noxref_28
cc_407 N_noxref_28_1 N_MM31_g 0.00165253f
cc_408 N_noxref_28_1 N_CLKB_13 0.000612844f
cc_409 N_noxref_28_1 N_NET0167_7 0.0360237f
cc_410 N_noxref_28_1 N_noxref_26_1 0.00769512f
cc_411 N_noxref_28_1 N_noxref_27_1 0.000469727f
x_PM_SDFLx2_ASAP7_75t_R%noxref_30 VSS N_noxref_30_1
+ PM_SDFLx2_ASAP7_75t_R%noxref_30
cc_412 N_noxref_30_1 N_CLKN_2 0.000184852f
cc_413 N_noxref_30_1 N_MM1_g 0.0107949f
cc_414 N_noxref_30_1 N_MM3_g 0.00149574f
cc_415 N_noxref_30_1 N_SI_1 0.00244743f
cc_416 N_noxref_30_1 N_PU1_2 0.00115942f
cc_417 N_noxref_30_1 N_PU1_10 0.0161892f
cc_418 N_noxref_30_1 N_PU1_9 0.0553171f
cc_419 N_noxref_30_1 N_NET0167_8 0.0371335f
x_PM_SDFLx2_ASAP7_75t_R%NET0167 VSS N_MM26_d N_MM5_s N_NET0167_7 N_NET0167_9
+ N_NET0167_1 N_NET0167_11 N_NET0167_12 N_NET0167_10 N_NET0167_8 N_NET0167_2
+ PM_SDFLx2_ASAP7_75t_R%NET0167
cc_420 N_NET0167_7 N_SE_1 0.00125998f
cc_421 N_NET0167_9 N_SE_10 0.000665382f
cc_422 N_NET0167_1 N_SE_8 0.000836735f
cc_423 N_NET0167_11 N_SE_7 0.00128214f
cc_424 N_NET0167_12 N_SE_10 0.0013577f
cc_425 N_NET0167_1 N_MM31_g 0.00158989f
cc_426 N_NET0167_11 N_SE_8 0.00388987f
cc_427 N_NET0167_10 N_SE_13 0.00440518f
cc_428 N_NET0167_7 N_MM31_g 0.0341766f
cc_429 N_NET0167_10 N_SEN_12 0.000325581f
cc_430 N_NET0167_10 N_SEN_16 0.000381233f
cc_431 N_NET0167_11 N_SEN_12 0.00109708f
cc_432 N_NET0167_10 N_SEN_14 0.00547666f
cc_433 N_NET0167_8 N_SI_1 0.00130032f
cc_434 N_NET0167_2 N_MM3_g 0.00153445f
cc_435 N_NET0167_8 N_MM3_g 0.0349042f
x_PM_SDFLx2_ASAP7_75t_R%PD1 VSS N_MM32_d N_MM5_d N_MM4_s N_PD1_8 N_PD1_2
+ N_PD1_9 N_PD1_7 N_PD1_1 PM_SDFLx2_ASAP7_75t_R%PD1
cc_436 N_PD1_8 N_CLKN_28 0.000153189f
cc_437 N_PD1_8 N_CLKN_2 0.0011149f
cc_438 N_PD1_2 N_MM1_g 0.0011671f
cc_439 N_PD1_9 N_CLKN_28 0.0023653f
cc_440 N_PD1_8 N_MM1_g 0.0355756f
cc_441 N_PD1_9 N_SE_13 0.00223299f
cc_442 N_PD1_9 N_MM27_g 0.000310135f
cc_443 N_PD1_9 N_SEN_12 0.000106357f
cc_444 N_PD1_9 N_SEN_14 0.000544416f
cc_445 N_PD1_9 N_SEN_16 0.00389418f
cc_446 N_PD1_7 N_D_1 0.000881293f
cc_447 N_PD1_1 N_MM30_g 0.00126331f
cc_448 N_PD1_9 N_D_5 0.00272066f
cc_449 N_PD1_7 N_MM30_g 0.0342671f
cc_450 N_PD1_9 N_SI_4 0.00043244f
cc_451 N_PD1_1 N_MM3_g 0.000757592f
cc_452 N_PD1_7 N_SI_1 0.000820741f
cc_453 N_PD1_9 N_SI_7 0.00251269f
cc_454 N_PD1_7 N_MM3_g 0.0334777f
cc_455 N_PD1_8 N_CLKB_1 0.000897958f
cc_456 N_PD1_9 N_CLKB_17 0.000742935f
cc_457 N_PD1_2 N_MM10_g 0.000866591f
cc_458 N_PD1_9 N_CLKB_22 0.000910038f
cc_459 N_PD1_8 N_MM10_g 0.0327525f
cc_460 N_PD1_8 N_MH_10 0.00114833f
cc_461 N_PD1_9 N_MH_15 0.000948957f
cc_462 N_PD1_2 N_MH_4 0.0036784f
cc_463 N_PD1_7 N_NET0167_10 0.00058352f
cc_464 N_PD1_9 N_NET0167_2 0.000634534f
cc_465 N_PD1_7 N_NET0167_8 0.000642602f
cc_466 N_PD1_1 N_NET0167_2 0.0038144f
cc_467 N_PD1_9 N_NET0167_10 0.00907615f
x_PM_SDFLx2_ASAP7_75t_R%SE VSS SE N_MM31_g N_MM0_g N_SE_9 N_SE_13 N_SE_8
+ N_SE_12 N_SE_1 N_SE_2 N_SE_10 N_SE_7 N_SE_11 PM_SDFLx2_ASAP7_75t_R%SE
x_PM_SDFLx2_ASAP7_75t_R%SEN VSS N_MM27_g N_MM0_d N_MM2_d N_SEN_3 N_SEN_4
+ N_SEN_13 N_SEN_14 N_SEN_1 N_SEN_15 N_SEN_11 N_SEN_10 N_SEN_12 N_SEN_16
+ PM_SDFLx2_ASAP7_75t_R%SEN
cc_468 N_SEN_3 N_SE_9 0.000160442f
cc_469 N_SEN_4 N_SE_9 0.000167851f
cc_470 N_SEN_13 N_SE_9 0.00803549f
cc_471 N_SEN_14 N_SE_13 0.000247294f
cc_472 N_SEN_1 N_SE_8 0.000309112f
cc_473 N_SEN_13 N_SE_12 0.000345458f
cc_474 N_SEN_15 N_SE_9 0.000409821f
cc_475 N_SEN_11 N_MM0_g 0.0159389f
cc_476 N_SEN_10 N_MM0_g 0.0536321f
cc_477 N_SEN_1 N_SE_1 0.00125681f
cc_478 N_SEN_12 N_SE_13 0.000479967f
cc_479 N_SEN_13 N_SE_13 0.000508708f
cc_480 N_SEN_4 N_SE_2 0.000685372f
cc_481 N_SEN_4 N_MM0_g 0.00133823f
cc_482 N_SEN_12 N_SE_8 0.00168423f
cc_483 N_SEN_3 N_MM0_g 0.00174322f
cc_484 N_SEN_11 N_SE_2 0.00174583f
cc_485 N_MM27_g N_MM31_g 0.00330887f
cc_486 N_SEN_16 N_SE_13 0.0649741f
*END of SDFLx2_ASAP7_75t_R.pxi
.ENDS
** Design:	SDFLx3_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "SDFLx3_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "SDFLx3_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_SDFLx3_ASAP7_75t_R%NET061 VSS 2 3 1
c1 1 VSS 0.000995471f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3780 $Y2=0.0675
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%noxref_33 VSS 1
c1 1 VSS 0.00447517f
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%noxref_34 VSS 1
c1 1 VSS 0.00479295f
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%noxref_35 VSS 1
c1 1 VSS 0.00541832f
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%noxref_31 VSS 1
c1 1 VSS 0.0034698f
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%noxref_32 VSS 1
c1 1 VSS 0.00368626f
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%noxref_36 VSS 1
c1 1 VSS 0.00535459f
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%QN VSS 32 24 25 35 42 43 45 13 19 3 15 4 18 1 2
+ 16 14
c1 1 VSS 0.0106725f
c2 2 VSS 0.0103505f
c3 3 VSS 0.00790815f
c4 4 VSS 0.00793668f
c5 13 VSS 0.00461845f
c6 14 VSS 0.00345898f
c7 15 VSS 0.00452949f
c8 16 VSS 0.00345357f
c9 17 VSS 0.0150294f
c10 18 VSS 0.0142594f
c11 19 VSS 0.00384414f
c12 20 VSS 0.00279929f
c13 21 VSS 0.00285596f
r1 16 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.3895 $Y=0.2025 $X2=1.4020 $Y2=0.2025
r2 45 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.3870 $Y=0.2025 $X2=1.3895 $Y2=0.2025
r3 43 41 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.3130 $Y=0.2025 $X2=1.3105 $Y2=0.2025
r4 2 41 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.2960 $Y=0.2025 $X2=1.3105 $Y2=0.2025
r5 15 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.2815 $Y=0.2025 $X2=1.2960 $Y2=0.2025
r6 42 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.2790 $Y=0.2025 $X2=1.2815 $Y2=0.2025
r7 4 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.4040 $Y=0.2025
+ $X2=1.4040 $Y2=0.2340
r8 2 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.2960 $Y=0.2025
+ $X2=1.2960 $Y2=0.2340
r9 38 39 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.4040
+ $Y=0.2340 $X2=1.4175 $Y2=0.2340
r10 37 38 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.3500
+ $Y=0.2340 $X2=1.4040 $Y2=0.2340
r11 36 37 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.2960
+ $Y=0.2340 $X2=1.3500 $Y2=0.2340
r12 18 36 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.2845
+ $Y=0.2340 $X2=1.2960 $Y2=0.2340
r13 21 33 0.624487 $w=2.20462e-08 $l=9.8e-09 $layer=M1 $thickness=3.6e-08
+ $X=1.4310 $Y=0.2340 $X2=1.4310 $Y2=0.2242
r14 21 39 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.4310 $Y=0.2340 $X2=1.4175 $Y2=0.2340
r15 14 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.3895 $Y=0.0675 $X2=1.4020 $Y2=0.0675
r16 35 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.3870 $Y=0.0675 $X2=1.3895 $Y2=0.0675
r17 32 33 0.291487 $w=1.3e-08 $l=1.2e-09 $layer=M1 $thickness=3.6e-08 $X=1.4310
+ $Y=0.2230 $X2=1.4310 $Y2=0.2242
r18 32 31 2.73998 $w=1.3e-08 $l=1.18e-08 $layer=M1 $thickness=3.6e-08 $X=1.4310
+ $Y=0.2230 $X2=1.4310 $Y2=0.2112
r19 30 31 15.4488 $w=1.3e-08 $l=6.62e-08 $layer=M1 $thickness=3.6e-08 $X=1.4310
+ $Y=0.1450 $X2=1.4310 $Y2=0.2112
r20 19 20 5.69636 $w=1.58e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.4310 $Y=0.0675 $X2=1.4310 $Y2=0.0360
r21 19 30 18.0722 $w=1.3e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=1.4310
+ $Y=0.0675 $X2=1.4310 $Y2=0.1450
r22 3 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.4040 $Y=0.0675
+ $X2=1.4040 $Y2=0.0360
r23 20 29 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.4310 $Y=0.0360 $X2=1.4175 $Y2=0.0360
r24 28 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.4040
+ $Y=0.0360 $X2=1.4175 $Y2=0.0360
r25 27 28 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.3500
+ $Y=0.0360 $X2=1.4040 $Y2=0.0360
r26 26 27 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.2960
+ $Y=0.0360 $X2=1.3500 $Y2=0.0360
r27 17 26 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.2845
+ $Y=0.0360 $X2=1.2960 $Y2=0.0360
r28 1 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.2960 $Y=0.0675
+ $X2=1.2960 $Y2=0.0360
r29 25 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.3130 $Y=0.0675 $X2=1.3105 $Y2=0.0675
r30 1 23 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.2960 $Y=0.0675 $X2=1.3105 $Y2=0.0675
r31 13 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.2815 $Y=0.0675 $X2=1.2960 $Y2=0.0675
r32 24 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.2790 $Y=0.0675 $X2=1.2815 $Y2=0.0675
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%D VSS 4 3 1 5
c1 1 VSS 0.00724305f
c2 3 VSS 0.0462133f
c3 4 VSS 0.00464529f
c4 5 VSS 0.0036858f
r1 5 7 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.1080 $X2=0.4050 $Y2=0.1215
r2 4 7 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1215
r3 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r4 4 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%NET062 VSS 14 27 7 9 1 11 12 10 8 2
c1 1 VSS 0.00639138f
c2 2 VSS 0.00558154f
c3 7 VSS 0.00468679f
c4 8 VSS 0.00322363f
c5 9 VSS 0.000875595f
c6 10 VSS 0.0175525f
c7 11 VSS 0.00131906f
c8 12 VSS 0.0020735f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0675 $X2=0.4840 $Y2=0.0675
r2 27 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4715 $Y2=0.0675
r3 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0675
+ $X2=0.4860 $Y2=0.0360
r4 23 24 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4475
+ $Y=0.0360 $X2=0.4860 $Y2=0.0360
r5 22 23 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4070
+ $Y=0.0360 $X2=0.4475 $Y2=0.0360
r6 21 22 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.3875
+ $Y=0.0360 $X2=0.4070 $Y2=0.0360
r7 20 21 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3605
+ $Y=0.0360 $X2=0.3875 $Y2=0.0360
r8 19 20 7.92845 $w=1.3e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3265
+ $Y=0.0360 $X2=0.3605 $Y2=0.0360
r9 10 12 1.03257 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3085 $Y=0.0360 $X2=0.2970 $Y2=0.0360
r10 10 19 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3085
+ $Y=0.0360 $X2=0.3265 $Y2=0.0360
r11 12 18 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.2970 $Y2=0.0540
r12 9 17 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0720 $X2=0.2970 $Y2=0.0900
r13 9 18 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0720 $X2=0.2970 $Y2=0.0540
r14 16 17 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2835 $Y=0.0900 $X2=0.2970 $Y2=0.0900
r15 11 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0900 $X2=0.2835 $Y2=0.0900
r16 11 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0900
+ $X2=0.2700 $Y2=0.0945
r17 1 15 23.8708 $w=2.02e-08 $l=4.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.2700 $Y=0.0540 $X2=0.2700 $Y2=0.0945
r18 14 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r19 7 13 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r20 1 7 1e-05
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%noxref_29 VSS 1
c1 1 VSS 0.00582495f
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%noxref_28 VSS 1
c1 1 VSS 0.00573324f
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%SE VSS 33 5 6 9 13 8 12 1 2 10 7 11
c1 1 VSS 0.00185567f
c2 2 VSS 0.00385954f
c3 5 VSS 0.0426614f
c4 6 VSS 0.0803916f
c5 7 VSS 0.00168936f
c6 8 VSS 0.000575907f
c7 9 VSS 0.00499659f
c8 10 VSS 0.00511274f
c9 11 VSS 0.00125994f
c10 12 VSS 0.00753306f
c11 13 VSS 0.0550085f
r1 1 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
r2 5 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r3 37 38 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2745
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r4 36 37 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2595
+ $Y=0.1350 $X2=0.2745 $Y2=0.1350
r5 35 36 0.699569 $w=1.3e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.1350 $X2=0.2595 $Y2=0.1350
r6 33 8 2.49951 $w=7.46154e-09 $l=1.95256e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.1340 $X2=0.2445 $Y2=0.1350
r7 8 35 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2445
+ $Y=0.1350 $X2=0.2565 $Y2=0.1350
r8 33 11 0.433689 $w=1.8e-08 $l=4.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.1340 $X2=0.2250 $Y2=0.1297
r9 11 31 3.53073 $w=1.4087e-08 $l=1.72e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.1297 $X2=0.2250 $Y2=0.1125
r10 10 27 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.2250 $Y=0.0360 $X2=0.2250
+ $Y2=0.0450
r11 30 31 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0900 $X2=0.2250 $Y2=0.1125
r12 29 30 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0675 $X2=0.2250 $Y2=0.0900
r13 7 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0495 $X2=0.2250 $Y2=0.0675
r14 7 27 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.2250 $Y=0.0495 $X2=0.2250
+ $Y2=0.0450
r15 7 10 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.0495 $X2=0.2250 $Y2=0.0360
r16 27 28 14.108 $w=1.3e-08 $l=6.05e-08 $layer=M2 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0450 $X2=0.2855 $Y2=0.0450
r17 25 28 109.716 $w=1.3e-08 $l=4.705e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.7560 $Y=0.0450 $X2=0.2855 $Y2=0.0450
r18 13 23 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=1.1905
+ $Y=0.0450 $X2=1.2150 $Y2=0.0450
r19 13 25 101.321 $w=1.3e-08 $l=4.345e-07 $layer=M2 $thickness=3.6e-08
+ $X=1.1905 $Y=0.0450 $X2=0.7560 $Y2=0.0450
r20 12 23 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=1.2150 $Y=0.0360 $X2=1.2150
+ $Y2=0.0450
r21 19 20 6.41272 $w=1.3e-08 $l=2.75e-08 $layer=M1 $thickness=3.6e-08 $X=1.2150
+ $Y=0.1085 $X2=1.2150 $Y2=0.1360
r22 18 19 8.51143 $w=1.3e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=1.2150
+ $Y=0.0720 $X2=1.2150 $Y2=0.1085
r23 9 18 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.2150
+ $Y=0.0495 $X2=1.2150 $Y2=0.0720
r24 9 12 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.2150 $Y=0.0495 $X2=1.2150 $Y2=0.0360
r25 9 23 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=1.2150 $Y=0.0495 $X2=1.2150
+ $Y2=0.0450
r26 17 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.2150 $Y=0.1380
+ $X2=1.2150 $Y2=0.1360
r27 6 2 1.49611 $w=1.91717e-07 $l=8e-09 $layer=LIG $thickness=5.46667e-08
+ $X=1.2150 $Y=0.1350 $X2=1.2150 $Y2=0.1270
r28 6 17 5.63117 $w=1.26721e-07 $l=3e-09 $layer=LIG $thickness=5.22105e-08
+ $X=1.2150 $Y=0.1350 $X2=1.2150 $Y2=0.1380
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%CLK VSS 11 3 4 6 1 5
c1 1 VSS 0.00307518f
c2 3 VSS 0.0599257f
c3 4 VSS 0.00149833f
c4 5 VSS 0.00465618f
c5 6 VSS 0.00196028f
r1 5 14 4.60559 $w=1.39091e-08 $l=2.74591e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0630 $X2=0.1030 $Y2=0.0900
r2 13 14 1.45753 $w=1.53529e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.0900 $X2=0.1030 $Y2=0.0900
r3 6 13 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0900 $X2=0.0945 $Y2=0.0900
r4 11 10 0.757867 $w=1.3e-08 $l=3.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1500 $X2=0.0810 $Y2=0.1467
r5 9 10 2.73998 $w=1.3e-08 $l=1.17e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1467
r6 8 9 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1235 $X2=0.0810 $Y2=0.1350
r7 4 8 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1100 $X2=0.0810 $Y2=0.1235
r8 4 6 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1100 $X2=0.0810 $Y2=0.0900
r9 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r10 1 9 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%NET063 VSS 12 13 27 28 9 7 1 2 8
c1 1 VSS 0.00533332f
c2 2 VSS 0.0053147f
c3 7 VSS 0.00333482f
c4 8 VSS 0.00335745f
c5 9 VSS 0.00273696f
r1 28 26 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r2 2 26 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r4 27 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r5 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4280 $Y2=0.1980
r6 21 22 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4185
+ $Y=0.1980 $X2=0.4280 $Y2=0.1980
r7 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1980 $X2=0.4185 $Y2=0.1980
r8 19 20 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.3875
+ $Y=0.1980 $X2=0.4050 $Y2=0.1980
r9 18 19 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3695
+ $Y=0.1980 $X2=0.3875 $Y2=0.1980
r10 17 18 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1980 $X2=0.3695 $Y2=0.1980
r11 16 17 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.1980 $X2=0.3510 $Y2=0.1980
r12 15 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1980 $X2=0.3375 $Y2=0.1980
r13 14 15 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3130
+ $Y=0.1980 $X2=0.3240 $Y2=0.1980
r14 9 14 0.699569 $w=1.3e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.3100
+ $Y=0.1980 $X2=0.3130 $Y2=0.1980
r15 1 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.1980
r16 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r17 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r18 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r19 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%SEN VSS 9 45 50 3 4 13 14 1 15 11 10 12 16
c1 1 VSS 0.0039046f
c2 3 VSS 0.00943925f
c3 4 VSS 0.00822429f
c4 9 VSS 0.0815967f
c5 10 VSS 0.00473746f
c6 11 VSS 0.00503622f
c7 12 VSS 0.00166699f
c8 13 VSS 0.00325061f
c9 14 VSS 0.000814545f
c10 15 VSS 0.00580974f
c11 16 VSS 0.0124058f
r1 50 49 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.2050 $Y=0.2025 $X2=1.2025 $Y2=0.2025
r2 11 49 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.1900 $Y=0.2025 $X2=1.2025 $Y2=0.2025
r3 4 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.1880 $Y=0.2295
+ $X2=1.1880 $Y2=0.2340
r4 45 44 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.2050 $Y=0.0675 $X2=1.2025 $Y2=0.0675
r5 10 44 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.1900 $Y=0.0675 $X2=1.2025 $Y2=0.0675
r6 41 42 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.1745
+ $Y=0.2340 $X2=1.1880 $Y2=0.2340
r7 15 37 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1610 $Y=0.2340 $X2=1.1610 $Y2=0.2125
r8 15 41 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1610 $Y=0.2340 $X2=1.1745 $Y2=0.2340
r9 3 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.1725 $Y=0.0405
+ $X2=1.1610 $Y2=0.0515
r10 3 10 4.30736 $w=5.12e-08 $l=2.95e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.1725 $Y=0.0405 $X2=1.1725 $Y2=0.0700
r11 36 37 15.7403 $w=1.3e-08 $l=6.75e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.1450 $X2=1.1610 $Y2=0.2125
r12 35 36 14.9241 $w=1.3e-08 $l=6.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0810 $X2=1.1610 $Y2=0.1450
r13 34 35 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0650 $X2=1.1610 $Y2=0.0810
r14 33 34 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0515 $X2=1.1610 $Y2=0.0650
r15 32 33 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0425 $X2=1.1610 $Y2=0.0515
r16 13 32 1.28254 $w=1.3e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0370 $X2=1.1610 $Y2=0.0425
r17 30 35 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=1.1610 $Y=0.0810
+ $X2=1.1610 $Y2=0.0810
r18 29 30 27.2832 $w=1.3e-08 $l=1.17e-07 $layer=M2 $thickness=3.6e-08 $X=1.0440
+ $Y=0.0810 $X2=1.1610 $Y2=0.0810
r19 28 29 29.3819 $w=1.3e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.9180
+ $Y=0.0810 $X2=1.0440 $Y2=0.0810
r20 27 28 67.1587 $w=1.3e-08 $l=2.88e-07 $layer=M2 $thickness=3.6e-08 $X=0.6300
+ $Y=0.0810 $X2=0.9180 $Y2=0.0810
r21 26 27 65.0599 $w=1.3e-08 $l=2.79e-07 $layer=M2 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0810 $X2=0.6300 $Y2=0.0810
r22 16 26 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.3395
+ $Y=0.0810 $X2=0.3510 $Y2=0.0810
r23 14 22 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.0720 $X2=0.3510 $Y2=0.0855
r24 14 26 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.3510 $Y=0.0720 $X2=0.3510
+ $Y2=0.0810
r25 22 23 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0855 $X2=0.3510 $Y2=0.0945
r26 22 26 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.3510 $Y=0.0855 $X2=0.3510
+ $Y2=0.0810
r27 21 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1080 $X2=0.3510 $Y2=0.0945
r28 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1215 $X2=0.3510 $Y2=0.1080
r29 12 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1215
r30 9 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r31 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
r32 4 11 1e-05
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%PD2 VSS 7 12 4 5 1
c1 1 VSS 0.00742561f
c2 4 VSS 0.00184273f
c3 5 VSS 0.00234046f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7040 $Y=0.2295 $X2=0.7165 $Y2=0.2295
r3 9 5 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.6765
+ $Y=0.2295 $X2=0.7020 $Y2=0.2295
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.6615
+ $Y=0.2295 $X2=0.6765 $Y2=0.2295
r5 1 8 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.6480
+ $Y=0.2295 $X2=0.6615 $Y2=0.2295
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.2295 $X2=0.6460 $Y2=0.2295
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.2295 $X2=0.6335 $Y2=0.2295
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%PD3 VSS 2 4 1
c1 1 VSS 0.0009112f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.0405 $X2=0.7065 $Y2=0.0405
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.0405 $X2=0.6895 $Y2=0.0405
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6895 $Y=0.0405 $X2=0.7065 $Y2=0.0405
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%PD5 VSS 7 12 1 5 4
c1 1 VSS 0.00742559f
c2 4 VSS 0.00187944f
c3 5 VSS 0.00237044f
r1 12 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9890 $Y=0.0405 $X2=0.9865 $Y2=0.0405
r2 5 11 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9740 $Y=0.0405 $X2=0.9865 $Y2=0.0405
r3 9 5 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.9585
+ $Y=0.0405 $X2=0.9720 $Y2=0.0405
r4 8 9 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.9435
+ $Y=0.0405 $X2=0.9585 $Y2=0.0405
r5 1 8 11.9937 $w=2.32e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08 $X=0.9180
+ $Y=0.0405 $X2=0.9435 $Y2=0.0405
r6 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9035 $Y=0.0405 $X2=0.9160 $Y2=0.0405
r7 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9010 $Y=0.0405 $X2=0.9035 $Y2=0.0405
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%SI VSS 14 3 5 6 7 1 4
c1 1 VSS 0.00578848f
c2 3 VSS 0.00731689f
c3 4 VSS 0.00310854f
c4 5 VSS 0.00300424f
c5 6 VSS 0.00356025f
c6 7 VSS 0.00369734f
r1 6 19 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1980 $X2=0.5130 $Y2=0.1765
r2 5 7 3.2503 $w=1.53684e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1540 $X2=0.5130 $Y2=0.1350
r3 5 19 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1540 $X2=0.5130 $Y2=0.1765
r4 7 16 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1350 $X2=0.4945 $Y2=0.1350
r5 15 16 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4845
+ $Y=0.1350 $X2=0.4945 $Y2=0.1350
r6 14 15 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4750
+ $Y=0.1350 $X2=0.4845 $Y2=0.1350
r7 14 4 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4750
+ $Y=0.1350 $X2=0.4635 $Y2=0.1350
r8 14 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4750 $Y=0.1350
+ $X2=0.4790 $Y2=0.1350
r9 11 12 4.43042 $w=1.53e-08 $l=7.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.4715
+ $Y=0.1350 $X2=0.4790 $Y2=0.1350
r10 9 11 1.86855 $w=1.78125e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.4675 $Y=0.1350 $X2=0.4715 $Y2=0.1350
r11 1 9 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.4575
+ $Y=0.1350 $X2=0.4675 $Y2=0.1350
r12 3 1 2.53453 $w=1.32811e-07 $l=1.5e-09 $layer=LIG $thickness=5.23243e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4575 $Y2=0.1350
r13 3 11 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4715 $Y2=0.1350
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%PD4 VSS 2 4 1
c1 1 VSS 0.00103f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9890 $Y=0.2295 $X2=0.9765 $Y2=0.2295
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9550 $Y=0.2295 $X2=0.9595 $Y2=0.2295
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9595 $Y=0.2295 $X2=0.9765 $Y2=0.2295
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%noxref_26 VSS 1
c1 1 VSS 0.00432558f
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%PU1 VSS 13 24 26 10 2 11 8 1 9
c1 1 VSS 0.00650224f
c2 2 VSS 0.00859741f
c3 8 VSS 0.00354215f
c4 9 VSS 0.0023747f
c5 10 VSS 0.00216315f
c6 11 VSS 0.0231093f
r1 26 25 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r2 10 25 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5420 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r3 9 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4840 $Y2=0.2025
r4 24 9 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r5 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5130 $Y=0.2025
+ $X2=0.4900 $Y2=0.2340
r6 20 21 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4810
+ $Y=0.2340 $X2=0.4900 $Y2=0.2340
r7 19 20 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4690
+ $Y=0.2340 $X2=0.4810 $Y2=0.2340
r8 18 19 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4540
+ $Y=0.2340 $X2=0.4690 $Y2=0.2340
r9 17 18 17.7224 $w=1.3e-08 $l=7.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.4540 $Y2=0.2340
r10 16 17 19.5879 $w=1.3e-08 $l=8.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2940
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r11 15 16 5.59655 $w=1.3e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.2940 $Y2=0.2340
r12 11 15 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2580
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r13 8 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2160
+ $X2=0.2700 $Y2=0.2340
r14 1 8 23.8708 $w=2.02e-08 $l=4.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.2700 $Y=0.1755 $X2=0.2700 $Y2=0.2160
r15 13 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r16 8 12 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r17 2 10 1e-05
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.00424559f
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%noxref_27 VSS 1
c1 1 VSS 0.00437026f
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%SS VSS 9 34 39 13 15 14 17 16 12 3 4 1 10 11
c1 1 VSS 0.00110935f
c2 3 VSS 0.0055653f
c3 4 VSS 0.00663772f
c4 9 VSS 0.0384164f
c5 10 VSS 0.00340948f
c6 11 VSS 0.00356123f
c7 12 VSS 0.00100091f
c8 13 VSS 0.00845562f
c9 14 VSS 0.00175941f
c10 15 VSS 0.00251702f
c11 16 VSS 0.00602217f
c12 17 VSS 0.00224388f
r1 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0655 $Y=0.2295 $X2=1.0780 $Y2=0.2295
r2 39 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0630 $Y=0.2295 $X2=1.0655 $Y2=0.2295
r3 4 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0800 $Y=0.2295
+ $X2=1.0800 $Y2=0.2340
r4 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.0800
+ $Y=0.2340 $X2=1.0935 $Y2=0.2340
r5 16 32 7.21452 $w=1.425e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.2340 $X2=1.1070 $Y2=0.1980
r6 16 37 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1070 $Y=0.2340 $X2=1.0935 $Y2=0.2340
r7 10 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.0655 $Y=0.0405 $X2=1.0780 $Y2=0.0405
r8 34 10 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.0630 $Y=0.0405 $X2=1.0655 $Y2=0.0405
r9 31 32 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.1440 $X2=1.1070 $Y2=0.1980
r10 14 30 8.95608 $w=1.36627e-08 $l=4.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1070 $Y=0.0810 $X2=1.1070 $Y2=0.0395
r11 14 31 14.691 $w=1.3e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.0810 $X2=1.1070 $Y2=0.1440
r12 3 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0800 $Y=0.0405
+ $X2=1.0800 $Y2=0.0360
r13 17 29 1.40651 $w=1.51875e-08 $l=1.45774e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.1070 $Y=0.0305 $X2=1.0935 $Y2=0.0360
r14 17 30 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.0305 $X2=1.1070 $Y2=0.0395
r15 28 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.0800
+ $Y=0.0360 $X2=1.0935 $Y2=0.0360
r16 27 28 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.0685
+ $Y=0.0360 $X2=1.0800 $Y2=0.0360
r17 26 27 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.0640
+ $Y=0.0360 $X2=1.0685 $Y2=0.0360
r18 25 26 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.0360 $X2=1.0640 $Y2=0.0360
r19 13 15 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0260 $Y=0.0360 $X2=0.9990 $Y2=0.0360
r20 13 25 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.0360 $X2=1.0530 $Y2=0.0360
r21 12 22 8.04505 $w=1.3e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.9990
+ $Y=0.0705 $X2=0.9990 $Y2=0.1050
r22 12 15 6.39593 $w=1.55565e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9990 $Y=0.0705 $X2=0.9990 $Y2=0.0360
r23 1 19 2.36633 $w=2.3e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.9990
+ $Y=0.1055 $X2=0.9990 $Y2=0.1055
r24 1 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.9990 $Y=0.1055
+ $X2=0.9990 $Y2=0.1050
r25 9 19 0.314665 $w=2.27e-07 $l=2.95e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.9990 $Y=0.1350 $X2=0.9990 $Y2=0.1055
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%MS VSS 10 43 46 50 52 3 15 13 12 1 17 11 4 18 19
+ 14 16
c1 1 VSS 0.00317647f
c2 3 VSS 0.00575065f
c3 4 VSS 0.00955879f
c4 10 VSS 0.0376965f
c5 11 VSS 0.003322f
c6 12 VSS 0.00315257f
c7 13 VSS 0.00266183f
c8 14 VSS 0.000856072f
c9 15 VSS 0.00355291f
c10 16 VSS 0.00188643f
c11 17 VSS 0.0011331f
c12 18 VSS 0.00136859f
c13 19 VSS 0.00117324f
c14 20 VSS 0.00294989f
r1 52 51 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8810 $Y=0.2295 $X2=0.8785 $Y2=0.2295
r2 13 51 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8660 $Y=0.2295 $X2=0.8785 $Y2=0.2295
r3 12 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.2295 $X2=0.8080 $Y2=0.2295
r4 50 12 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.2295 $X2=0.7955 $Y2=0.2295
r5 47 13 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8370 $Y=0.2295 $X2=0.8640 $Y2=0.2295
r6 4 47 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08 $X=0.8100
+ $Y=0.2295 $X2=0.8370 $Y2=0.2295
r7 4 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8100 $Y=0.2295
+ $X2=0.8100 $Y2=0.2340
r8 15 20 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.2340 $X2=0.8370 $Y2=0.2340
r9 46 45 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8270 $Y=0.0405 $X2=0.8245 $Y2=0.0405
r10 44 45 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8200 $Y=0.0405 $X2=0.8245 $Y2=0.0405
r11 3 44 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8080 $Y=0.0405 $X2=0.8200 $Y2=0.0405
r12 11 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.0405 $X2=0.8080 $Y2=0.0405
r13 43 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.0405 $X2=0.7955 $Y2=0.0405
r14 20 39 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.2340 $X2=0.8370 $Y2=0.2160
r15 3 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8100 $Y=0.0405
+ $X2=0.8100 $Y2=0.0535
r16 38 39 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1870 $X2=0.8370 $Y2=0.2160
r17 37 38 4.89699 $w=1.3e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1660 $X2=0.8370 $Y2=0.1870
r18 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1525 $X2=0.8370 $Y2=0.1660
r19 35 36 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1310 $X2=0.8370 $Y2=0.1525
r20 34 35 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1115 $X2=0.8370 $Y2=0.1310
r21 17 31 1.15159 $w=1.75e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1000 $X2=0.8370 $Y2=0.0900
r22 17 34 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1000 $X2=0.8370 $Y2=0.1115
r23 16 32 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0625 $X2=0.8100 $Y2=0.0720
r24 16 33 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0625 $X2=0.8100 $Y2=0.0535
r25 30 31 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8235 $Y=0.0900 $X2=0.8370 $Y2=0.0900
r26 19 28 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.0900 $X2=0.7965 $Y2=0.0900
r27 19 30 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.0900 $X2=0.8235 $Y2=0.0900
r28 19 32 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0900 $X2=0.8100 $Y2=0.0720
r29 27 28 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.7740
+ $Y=0.0900 $X2=0.7965 $Y2=0.0900
r30 14 27 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7470
+ $Y=0.0900 $X2=0.7740 $Y2=0.0900
r31 14 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7470 $Y=0.0900
+ $X2=0.7500 $Y2=0.0900
r32 14 18 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7470
+ $Y=0.0900 $X2=0.7290 $Y2=0.0900
r33 25 26 5.02115 $w=1.53e-08 $l=8.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.7415 $Y=0.0900 $X2=0.7500 $Y2=0.0900
r34 23 25 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.7385 $Y=0.0900 $X2=0.7415 $Y2=0.0900
r35 1 23 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.7285
+ $Y=0.0900 $X2=0.7385 $Y2=0.0900
r36 1 22 2.48102 $w=2.2e-08 $l=5e-10 $layer=LIG $thickness=4.8e-08 $X=0.7285
+ $Y=0.0900 $X2=0.7290 $Y2=0.0900
r37 22 25 1.47681 $w=1.53e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7290 $Y=0.0900 $X2=0.7415 $Y2=0.0900
r38 10 22 0.314665 $w=2.27e-07 $l=4.5e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.7290 $Y=0.1350 $X2=0.7290 $Y2=0.0900
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%PD1 VSS 12 13 29 8 2 9 7 1
c1 1 VSS 0.00350932f
c2 2 VSS 0.00380949f
c3 7 VSS 0.00294155f
c4 8 VSS 0.0022742f
c5 9 VSS 0.00243992f
r1 29 28 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.0675 $X2=0.6085 $Y2=0.0675
r2 27 28 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6040 $Y=0.0675 $X2=0.6085 $Y2=0.0675
r3 8 27 0.123457 $w=8.1e-08 $l=1e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.0675 $X2=0.6040 $Y2=0.0675
r4 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0675
+ $X2=0.5900 $Y2=0.0720
r5 23 24 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.5805
+ $Y=0.0720 $X2=0.5900 $Y2=0.0720
r6 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0720 $X2=0.5805 $Y2=0.0720
r7 21 22 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.0720 $X2=0.5670 $Y2=0.0720
r8 20 21 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0720 $X2=0.5400 $Y2=0.0720
r9 19 20 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5020
+ $Y=0.0720 $X2=0.5130 $Y2=0.0720
r10 18 19 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4805
+ $Y=0.0720 $X2=0.5020 $Y2=0.0720
r11 17 18 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.4540
+ $Y=0.0720 $X2=0.4805 $Y2=0.0720
r12 16 17 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4440
+ $Y=0.0720 $X2=0.4540 $Y2=0.0720
r13 15 16 1.63233 $w=1.3e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.4370
+ $Y=0.0720 $X2=0.4440 $Y2=0.0720
r14 14 15 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4280
+ $Y=0.0720 $X2=0.4370 $Y2=0.0720
r15 9 14 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4205
+ $Y=0.0720 $X2=0.4280 $Y2=0.0720
r16 1 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4280 $Y2=0.0720
r17 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r18 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r19 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0675 $X2=0.4320 $Y2=0.0675
r20 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4175 $Y2=0.0675
r21 2 8 1e-05
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.00423343f
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%noxref_30 VSS 1
c1 1 VSS 0.0124552f
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%MH VSS 9 55 59 62 66 10 3 21 17 1 4 12 14 18 20
+ 16 19 15
c1 1 VSS 0.000217469f
c2 3 VSS 0.00473518f
c3 4 VSS 0.00495888f
c4 9 VSS 0.036124f
c5 10 VSS 0.00226938f
c6 11 VSS 9.97604e-20
c7 12 VSS 0.00211058f
c8 13 VSS 6.70519e-20
c9 14 VSS 0.00910063f
c10 15 VSS 0.00778544f
c11 16 VSS 0.00174644f
c12 17 VSS 0.000617839f
c13 18 VSS 0.000950246f
c14 19 VSS 0.00298446f
c15 20 VSS 5.93462e-20
c16 21 VSS 0.00268982f
r1 66 65 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.2295 $X2=0.6085 $Y2=0.2295
r2 64 65 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6040 $Y=0.2295 $X2=0.6085 $Y2=0.2295
r3 3 64 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5920 $Y=0.2295 $X2=0.6040 $Y2=0.2295
r4 13 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2295 $X2=0.5920 $Y2=0.2295
r5 60 61 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.1890 $X2=0.5840 $Y2=0.1890
r6 62 60 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.1890 $X2=0.5795 $Y2=0.1890
r7 12 61 0.185185 $w=5.4e-08 $l=1e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.1890 $X2=0.5840 $Y2=0.1890
r8 12 3 0.518519 $w=3.9e-08 $l=4.05494e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.1890 $X2=0.5920 $Y2=0.2295
r9 59 58 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r10 57 58 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6580 $Y=0.0405 $X2=0.6625 $Y2=0.0405
r11 4 57 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6460 $Y=0.0405 $X2=0.6580 $Y2=0.0405
r12 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0405 $X2=0.6460 $Y2=0.0405
r13 10 4 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0810 $X2=0.6460 $Y2=0.0810
r14 55 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.0810 $X2=0.6335 $Y2=0.0810
r15 3 47 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2295
+ $X2=0.5900 $Y2=0.2340
r16 4 41 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.0405
+ $X2=0.6440 $Y2=0.0360
r17 44 45 1.63233 $w=1.3e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.5990
+ $Y=0.2340 $X2=0.6060 $Y2=0.2340
r18 44 47 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5990
+ $Y=0.2340 $X2=0.5900 $Y2=0.2340
r19 43 45 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.6105
+ $Y=0.2340 $X2=0.6060 $Y2=0.2340
r20 42 43 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6305
+ $Y=0.2340 $X2=0.6105 $Y2=0.2340
r21 14 21 4.53042 $w=1.46981e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6665 $Y=0.2340 $X2=0.6930 $Y2=0.2340
r22 14 42 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.6665
+ $Y=0.2340 $X2=0.6305 $Y2=0.2340
r23 15 39 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.6530
+ $Y=0.0360 $X2=0.6705 $Y2=0.0360
r24 15 41 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6530
+ $Y=0.0360 $X2=0.6440 $Y2=0.0360
r25 21 38 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.2340 $X2=0.6930 $Y2=0.2160
r26 19 33 2.43171 $w=1.804e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6930 $Y=0.0360 $X2=0.6930 $Y2=0.0535
r27 19 39 3.59766 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.0360 $X2=0.6705 $Y2=0.0360
r28 37 38 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1980 $X2=0.6930 $Y2=0.2160
r29 36 37 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1800 $X2=0.6930 $Y2=0.1980
r30 35 36 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1680 $X2=0.6930 $Y2=0.1800
r31 34 35 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1590 $X2=0.6930 $Y2=0.1680
r32 17 20 2.43413 $w=1.59032e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6930 $Y=0.1465 $X2=0.6930 $Y2=0.1310
r33 17 34 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1465 $X2=0.6930 $Y2=0.1590
r34 32 33 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.0625 $X2=0.6930 $Y2=0.0535
r35 31 32 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.0720 $X2=0.6930 $Y2=0.0625
r36 30 31 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.0900 $X2=0.6930 $Y2=0.0720
r37 29 30 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1025 $X2=0.6930 $Y2=0.0900
r38 16 20 2.78392 $w=1.56471e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6930 $Y=0.1140 $X2=0.6930 $Y2=0.1310
r39 16 29 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1140 $X2=0.6930 $Y2=0.1025
r40 20 28 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1310 $X2=0.7110 $Y2=0.1310
r41 27 28 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1310 $X2=0.7110 $Y2=0.1310
r42 18 26 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.1310 $X2=0.7830 $Y2=0.1310
r43 18 27 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.1310 $X2=0.7290 $Y2=0.1310
r44 1 23 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.7830
+ $Y=0.1310 $X2=0.7830 $Y2=0.1310
r45 1 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7830 $Y=0.1310
+ $X2=0.7830 $Y2=0.1310
r46 9 23 0.314665 $w=2.27e-07 $l=4e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.7830 $Y=0.1350 $X2=0.7830 $Y2=0.1310
r47 3 12 1e-05
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%CLKB VSS 11 12 61 63 13 22 16 5 19 15 6 20 14 17
+ 18 2 1 21
c1 1 VSS 0.000148262f
c2 2 VSS 0.000213148f
c3 5 VSS 0.00733852f
c4 6 VSS 0.00724018f
c5 11 VSS 0.0044918f
c6 12 VSS 0.00460296f
c7 13 VSS 0.00745879f
c8 14 VSS 0.00750874f
c9 15 VSS 0.00646166f
c10 16 VSS 0.00361469f
c11 17 VSS 0.000128357f
c12 18 VSS 0.000485179f
c13 19 VSS 0.00590553f
c14 20 VSS 0.00306033f
c15 21 VSS 0.000164032f
c16 22 VSS 0.0197055f
r1 14 6 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1600 $Y2=0.2160
r2 63 14 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r3 6 56 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r4 13 5 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1600 $Y2=0.0540
r5 61 13 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r6 56 57 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r7 15 56 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1505
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r8 5 53 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r9 20 49 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.1890 $Y2=0.2160
r10 20 57 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2340 $X2=0.1755 $Y2=0.2340
r11 53 54 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r12 19 44 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1890 $Y2=0.0630
r13 19 54 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1755 $Y2=0.0360
r14 1 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6210 $Y=0.1350
+ $X2=0.6210 $Y2=0.1395
r15 11 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1350
r16 48 49 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1980 $X2=0.1890 $Y2=0.2160
r17 47 48 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1765 $X2=0.1890 $Y2=0.1980
r18 46 47 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1630 $X2=0.1890 $Y2=0.1765
r19 45 46 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1530 $X2=0.1890 $Y2=0.1630
r20 43 44 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0900 $X2=0.1890 $Y2=0.0630
r21 42 43 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1100 $X2=0.1890 $Y2=0.0900
r22 16 42 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1325 $X2=0.1890 $Y2=0.1100
r23 16 45 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1325 $X2=0.1890 $Y2=0.1530
r24 21 39 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1620 $X2=0.6210 $Y2=0.1395
r25 21 33 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.6210 $Y=0.1620 $X2=0.6210
+ $Y2=0.1530
r26 17 39 5.47996 $w=1.3e-08 $l=2.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1160 $X2=0.6210 $Y2=0.1395
r27 37 38 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1530 $X2=0.2045 $Y2=0.1530
r28 37 45 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1890 $Y=0.1530
+ $X2=0.1890 $Y2=0.1530
r29 35 38 16.2067 $w=1.3e-08 $l=6.95e-08 $layer=M2 $thickness=3.6e-08 $X=0.2740
+ $Y=0.1530 $X2=0.2045 $Y2=0.1530
r30 33 34 15.2739 $w=1.3e-08 $l=6.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1530 $X2=0.6865 $Y2=0.1530
r31 33 39 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.6210 $Y=0.1530 $X2=0.6210
+ $Y2=0.1395
r32 32 33 34.1623 $w=1.3e-08 $l=1.465e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.4745 $Y=0.1530 $X2=0.6210 $Y2=0.1530
r33 32 35 46.7545 $w=1.3e-08 $l=2.005e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.4745 $Y=0.1530 $X2=0.2740 $Y2=0.1530
r34 22 31 18.3054 $w=1.3e-08 $l=7.85e-08 $layer=M2 $thickness=3.6e-08 $X=0.8125
+ $Y=0.1530 $X2=0.8910 $Y2=0.1530
r35 22 34 29.3819 $w=1.3e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.8125
+ $Y=0.1530 $X2=0.6865 $Y2=0.1530
r36 29 31 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.8910 $Y=0.1440
+ $X2=0.8910 $Y2=0.1530
r37 18 29 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1135 $X2=0.8910 $Y2=0.1440
r38 12 2 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.8910
+ $Y=0.1350 $X2=0.8910 $Y2=0.1350
r39 2 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8910 $Y=0.1350
+ $X2=0.8910 $Y2=0.1440
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%CLKN VSS 16 17 18 19 20 101 103 30 27 26 31 8 22
+ 21 33 9 1 35 25 23 2 28 34 10 5 29 3 32 24
c1 1 VSS 0.00150493f
c2 2 VSS 0.000252245f
c3 3 VSS 5.46221e-20
c4 4 VSS 1e-36
c5 5 VSS 0.000273532f
c6 8 VSS 0.00776474f
c7 9 VSS 0.00800184f
c8 10 VSS 0.00382808f
c9 16 VSS 0.0593152f
c10 17 VSS 0.00580365f
c11 18 VSS 0.00508225f
c12 19 VSS 0.00437088f
c13 20 VSS 0.00534604f
c14 21 VSS 0.00646115f
c15 22 VSS 0.00638007f
c16 23 VSS 0.00788445f
c17 24 VSS 0.0017795f
c18 25 VSS 0.00463367f
c19 26 VSS 0.00375908f
c20 27 VSS 0.00114558f
c21 28 VSS 0.0025362f
c22 29 VSS 0.00137914f
c23 30 VSS 0.00366487f
c24 31 VSS 0.00197507f
c25 32 VSS 0.00396616f
c26 33 VSS 0.00138132f
c27 34 VSS 0.000588057f
c28 35 VSS 0.0299541f
r1 103 102 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r2 22 102 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r3 101 100 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r4 21 100 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r5 9 98 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0550 $Y2=0.2340
r6 8 95 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0550 $Y2=0.0360
r7 97 98 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.2340 $X2=0.0550 $Y2=0.2340
r8 26 97 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0460 $Y2=0.2340
r9 26 32 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0180 $Y2=0.2340
r10 94 95 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.0360 $X2=0.0550 $Y2=0.0360
r11 25 94 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0460 $Y2=0.0360
r12 25 30 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0180 $Y2=0.0360
r13 32 92 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.2340 $X2=0.0180 $Y2=0.2160
r14 30 91 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.0360 $X2=0.0180 $Y2=0.0630
r15 1 83 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
r16 16 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r17 24 31 1.81469 $w=1.6125e-08 $l=1.35831e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.2025 $X2=0.0165 $Y2=0.1890
r18 24 92 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.2025 $X2=0.0180 $Y2=0.2160
r19 90 91 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0900 $X2=0.0180 $Y2=0.0630
r20 89 90 9.67737 $w=1.3e-08 $l=4.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1315 $X2=0.0180 $Y2=0.0900
r21 23 31 2.63085 $w=1.54194e-08 $l=1.7066e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1720 $X2=0.0165 $Y2=0.1890
r22 23 89 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1720 $X2=0.0180 $Y2=0.1315
r23 2 74 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1355
+ $X2=0.5670 $Y2=0.1350
r24 17 2 3.19489 $w=1.24e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1355
r25 33 69 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.1350 $Y=0.1980 $X2=0.1350
+ $Y2=0.1890
r26 83 84 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1540
r27 81 84 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1720 $X2=0.1350 $Y2=0.1540
r28 27 69 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.1350 $Y=0.1845 $X2=0.1350
+ $Y2=0.1890
r29 27 81 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1845 $X2=0.1350 $Y2=0.1720
r30 27 33 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1845 $X2=0.1350 $Y2=0.1980
r31 78 79 1.90199 $w=1.38333e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.0255 $Y=0.1890 $X2=0.0345 $Y2=0.1890
r32 31 78 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0165
+ $Y=0.1890 $X2=0.0255 $Y2=0.1890
r33 34 71 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.1980 $X2=0.5670 $Y2=0.1845
r34 34 62 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.5670 $Y=0.1980 $X2=0.5670
+ $Y2=0.1890
r35 74 75 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1485
r36 72 75 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1620 $X2=0.5670 $Y2=0.1485
r37 28 71 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1755 $X2=0.5670 $Y2=0.1845
r38 28 72 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1755 $X2=0.5670 $Y2=0.1620
r39 69 70 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1890 $X2=0.1595 $Y2=0.1890
r40 68 69 11.8927 $w=1.3e-08 $l=5.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.0840
+ $Y=0.1890 $X2=0.1350 $Y2=0.1890
r41 67 68 11.8927 $w=1.3e-08 $l=5.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.0330
+ $Y=0.1890 $X2=0.0840 $Y2=0.1890
r42 67 79 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.0330 $Y=0.1890
+ $X2=0.0345 $Y2=0.1890
r43 63 64 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.6480
+ $Y=0.1890 $X2=0.7290 $Y2=0.1890
r44 62 63 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1890 $X2=0.6480 $Y2=0.1890
r45 62 71 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.5670 $Y=0.1890 $X2=0.5670
+ $Y2=0.1845
r46 35 62 46.7546 $w=1.3e-08 $l=2.005e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.3665 $Y=0.1890 $X2=0.5670 $Y2=0.1890
r47 35 70 48.2703 $w=1.3e-08 $l=2.07e-07 $layer=M2 $thickness=3.6e-08 $X=0.3665
+ $Y=0.1890 $X2=0.1595 $Y2=0.1890
r48 5 59 2.78395 $w=2.4e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.9450
+ $Y=0.1780 $X2=0.9450 $Y2=0.1780
r49 20 5 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.9450 $Y=0.1350 $X2=0.9450 $Y2=0.1780
r50 3 52 2.78395 $w=2.4e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.6750
+ $Y=0.1780 $X2=0.6750 $Y2=0.1780
r51 18 3 3.09861 $w=1.12261e-07 $l=4.3e-08 $layer=LIG $thickness=5.14783e-08
+ $X=0.6750 $Y=0.1350 $X2=0.6750 $Y2=0.1780
r52 60 64 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.7290 $Y=0.1845
+ $X2=0.7290 $Y2=0.1890
r53 29 60 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1680 $X2=0.7290 $Y2=0.1845
r54 58 59 6.83711 $w=2.22e-08 $l=1.5e-09 $layer=LISD $thickness=2.7e-08
+ $X=0.9435 $Y=0.1780 $X2=0.9450 $Y2=0.1780
r55 57 58 12.9145 $w=2.22e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9180 $Y=0.1780 $X2=0.9435 $Y2=0.1780
r56 56 57 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9045 $Y=0.1780 $X2=0.9180 $Y2=0.1780
r57 55 56 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8910 $Y=0.1780 $X2=0.9045 $Y2=0.1780
r58 54 55 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8775 $Y=0.1780 $X2=0.8910 $Y2=0.1780
r59 53 54 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8640 $Y=0.1780 $X2=0.8775 $Y2=0.1780
r60 51 52 12.9145 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6885 $Y=0.1780 $X2=0.6750 $Y2=0.1780
r61 50 51 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7155 $Y=0.1780 $X2=0.6885 $Y2=0.1780
r62 48 49 6.07743 $w=2.22e-08 $l=1.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7290 $Y=0.1780 $X2=0.7410 $Y2=0.1780
r63 48 60 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7290 $Y=0.1780
+ $X2=0.7290 $Y2=0.1845
r64 47 48 5.31775 $w=2.22e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7185 $Y=0.1780 $X2=0.7290 $Y2=0.1780
r65 47 50 1.51936 $w=2.22e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.7185
+ $Y=0.1780 $X2=0.7155 $Y2=0.1780
r66 46 49 4.55807 $w=2.22e-08 $l=9e-09 $layer=LISD $thickness=2.7e-08 $X=0.7500
+ $Y=0.1780 $X2=0.7410 $Y2=0.1780
r67 45 46 6.07743 $w=2.22e-08 $l=1.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7620 $Y=0.1780 $X2=0.7500 $Y2=0.1780
r68 44 45 4.05162 $w=2.22e-08 $l=8e-09 $layer=LISD $thickness=2.7e-08 $X=0.7700
+ $Y=0.1780 $X2=0.7620 $Y2=0.1780
r69 43 44 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7835 $Y=0.1780 $X2=0.7700 $Y2=0.1780
r70 42 43 6.58388 $w=2.22e-08 $l=1.3e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7965 $Y=0.1780 $X2=0.7835 $Y2=0.1780
r71 41 42 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8100 $Y=0.1780 $X2=0.7965 $Y2=0.1780
r72 10 41 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8370 $Y=0.1780 $X2=0.8100 $Y2=0.1780
r73 10 53 13.6742 $w=2.22e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8370 $Y=0.1780 $X2=0.8640 $Y2=0.1780
r74 4 40 2.78395 $w=2.4e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.8370
+ $Y=0.1780 $X2=0.8370 $Y2=0.1780
r75 4 10 10.3807 $w=2.30357e-08 $l=0 $layer=LISD $thickness=3.675e-08 $X=0.8370
+ $Y=0.1780 $X2=0.8370 $Y2=0.1780
r76 19 40 0.314665 $w=2.27e-07 $l=4.3e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.8370 $Y=0.1350 $X2=0.8370 $Y2=0.1780
r77 9 22 1e-05
r78 8 21 1e-05
.ends

.subckt PM_SDFLx3_ASAP7_75t_R%SH VSS 11 12 13 14 83 86 88 91 16 17 23 25 15 6
+ 20 18 19 5 22 24 2 27 1 21 26
c1 1 VSS 0.0024806f
c2 2 VSS 0.0148123f
c3 5 VSS 0.00684057f
c4 6 VSS 0.00697309f
c5 11 VSS 0.0386518f
c6 12 VSS 0.0815734f
c7 13 VSS 0.081305f
c8 14 VSS 0.0809895f
c9 15 VSS 0.00494786f
c10 16 VSS 0.00515575f
c11 17 VSS 0.00889377f
c12 18 VSS 0.00247168f
c13 19 VSS 0.00213443f
c14 20 VSS 0.00208334f
c15 21 VSS 0.00106037f
c16 22 VSS 0.00501557f
c17 23 VSS 0.00726265f
c18 24 VSS 0.00306646f
c19 25 VSS 0.000990843f
c20 26 VSS 0.00121664f
c21 27 VSS 0.00479268f
r1 91 90 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8810 $Y=0.0405 $X2=0.8785 $Y2=0.0405
r2 5 90 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8660 $Y=0.0405 $X2=0.8785 $Y2=0.0405
r3 87 5 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8540 $Y=0.0405 $X2=0.8660 $Y2=0.0405
r4 15 87 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.0405 $X2=0.8540 $Y2=0.0405
r5 88 15 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.0405 $X2=0.8495 $Y2=0.0405
r6 86 85 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9350 $Y=0.2295 $X2=0.9325 $Y2=0.2295
r7 84 85 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9280 $Y=0.2295 $X2=0.9325 $Y2=0.2295
r8 6 84 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9160 $Y=0.2295 $X2=0.9280 $Y2=0.2295
r9 16 6 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9035 $Y=0.2295 $X2=0.9160 $Y2=0.2295
r10 83 16 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9010 $Y=0.2295 $X2=0.9035 $Y2=0.2295
r11 14 75 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=1.3770
+ $Y=0.1350 $X2=1.3770 $Y2=0.1360
r12 13 69 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=1.3230
+ $Y=0.1350 $X2=1.3230 $Y2=0.1360
r13 12 61 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=1.2690 $Y=0.1350 $X2=1.2690 $Y2=0.1360
r14 5 59 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.0405
+ $X2=0.8640 $Y2=0.0360
r15 6 54 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.9180 $Y=0.2295
+ $X2=0.9180 $Y2=0.2340
r16 73 75 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.3645 $Y=0.1360 $X2=1.3770 $Y2=0.1360
r17 72 73 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.3500 $Y=0.1360 $X2=1.3645 $Y2=0.1360
r18 70 72 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.3355 $Y=0.1360 $X2=1.3500 $Y2=0.1360
r19 69 70 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.3230 $Y=0.1360 $X2=1.3355 $Y2=0.1360
r20 67 69 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.3105 $Y=0.1360 $X2=1.3230 $Y2=0.1360
r21 66 67 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.2960 $Y=0.1360 $X2=1.3105 $Y2=0.1360
r22 64 66 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.2815 $Y=0.1360 $X2=1.2960 $Y2=0.1360
r23 62 64 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=1.2785 $Y=0.1360 $X2=1.2815 $Y2=0.1360
r24 61 62 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=1.2690
+ $Y=0.1360 $X2=1.2785 $Y2=0.1360
r25 2 61 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=1.2595
+ $Y=0.1360 $X2=1.2690 $Y2=0.1360
r26 59 60 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.0360 $X2=0.8775 $Y2=0.0360
r27 57 60 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.0360 $X2=0.8775 $Y2=0.0360
r28 56 57 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.9020
+ $Y=0.0360 $X2=0.8910 $Y2=0.0360
r29 17 24 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.9200
+ $Y=0.0360 $X2=0.9450 $Y2=0.0360
r30 17 56 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.9200
+ $Y=0.0360 $X2=0.9020 $Y2=0.0360
r31 54 55 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.2340 $X2=0.9315 $Y2=0.2340
r32 23 55 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.2340 $X2=0.9315 $Y2=0.2340
r33 51 61 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.2690 $Y=0.1445
+ $X2=1.2690 $Y2=0.1360
r34 22 51 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.2690
+ $Y=0.1085 $X2=1.2690 $Y2=0.1445
r35 24 45 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.0360 $X2=0.9450 $Y2=0.0630
r36 19 40 6.50021 $w=1.33448e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.1980 $X2=0.9450 $Y2=0.1690
r37 19 23 7.21452 $w=1.425e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.1980 $X2=0.9450 $Y2=0.2340
r38 49 51 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=1.2690 $Y=0.1530
+ $X2=1.2690 $Y2=0.1445
r39 48 49 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=1.2445
+ $Y=0.1530 $X2=1.2690 $Y2=0.1530
r40 47 48 9.91056 $w=1.3e-08 $l=4.25e-08 $layer=M2 $thickness=3.6e-08 $X=1.2020
+ $Y=0.1530 $X2=1.2445 $Y2=0.1530
r41 46 47 32.0636 $w=1.3e-08 $l=1.375e-07 $layer=M2 $thickness=3.6e-08
+ $X=1.0645 $Y=0.1530 $X2=1.2020 $Y2=0.1530
r42 27 46 27.8662 $w=1.3e-08 $l=1.195e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.9450 $Y=0.1530 $X2=1.0645 $Y2=0.1530
r43 27 41 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.9450 $Y=0.1530 $X2=0.9450
+ $Y2=0.1485
r44 44 45 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.0900 $X2=0.9450 $Y2=0.0630
r45 43 44 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1000 $X2=0.9450 $Y2=0.0900
r46 42 43 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1100 $X2=0.9450 $Y2=0.1000
r47 18 41 3.96423 $w=1.3e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1315 $X2=0.9450 $Y2=0.1485
r48 18 42 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1315 $X2=0.9450 $Y2=0.1100
r49 39 40 0.4592 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1645 $X2=0.9450 $Y2=0.1690
r50 25 39 0.714311 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1575 $X2=0.9450 $Y2=0.1645
r51 25 41 1.50855 $w=1.55e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1575 $X2=0.9450 $Y2=0.1485
r52 25 27 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.9450 $Y=0.1575 $X2=0.9450
+ $Y2=0.1530
r53 38 40 4.4015 $w=1.35e-08 $l=2.78927e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9720 $Y=0.1620 $X2=0.9450 $Y2=0.1690
r54 37 38 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9990
+ $Y=0.1620 $X2=0.9720 $Y2=0.1620
r55 20 26 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0260 $Y=0.1620 $X2=1.0530 $Y2=0.1620
r56 20 37 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.1620 $X2=0.9990 $Y2=0.1620
r57 26 35 0.915974 $w=2.10182e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0530 $Y=0.1620 $X2=1.0530 $Y2=0.1510
r58 34 35 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1400 $X2=1.0530 $Y2=0.1510
r59 21 34 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1250 $X2=1.0530 $Y2=0.1400
r60 1 31 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=1.0530
+ $Y=0.1400 $X2=1.0530 $Y2=0.1400
r61 1 34 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.0530 $Y=0.1400
+ $X2=1.0530 $Y2=0.1400
r62 11 31 0.314665 $w=2.27e-07 $l=5e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.0530 $Y=0.1350 $X2=1.0530 $Y2=0.1400
.ends


*
.SUBCKT SDFLx3_ASAP7_75t_R VSS VDD CLK SE D SI QN
*
* VSS VSS
* VDD VDD
* CLK CLK
* SE SE
* D D
* SI SI
* QN QN
*
*

MM20 N_MM20_d N_MM20_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM23 N_MM23_d N_MM22_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM26 N_MM26_d N_MM31_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM29 N_MM29_d N_MM27_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM32 N_MM32_d N_MM30_g N_MM32_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM3_g N_MM5_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM10_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM6 N_MM6_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM12 N_MM12_d N_MM12_g N_MM12_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM17 N_MM17_d N_MM17_g N_MM17_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM16 N_MM16_d N_MM16_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM14 N_MM14_d N_MM14_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM0 N_MM0_d N_MM0_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24 N_MM24_d N_MM24_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@3 N_MM24@3_d N_MM24@3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@2 N_MM24@2_d N_MM24@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM21 N_MM21_d N_MM20_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM22 N_MM22_d N_MM22_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM31 N_MM31_d N_MM31_g N_MM31_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM27 N_MM27_d N_MM27_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM30 N_MM30_d N_MM30_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g N_MM3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM13 N_MM13_d N_MM17_g N_MM13_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM18 N_MM18_d N_MM18_g N_MM18_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM19 N_MM19_d N_MM16_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM15 N_MM15_d N_MM14_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM2 N_MM2_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25 N_MM25_d N_MM24_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@3 N_MM25@3_d N_MM24@3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@2 N_MM25@2_d N_MM24@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "SDFLx3_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "SDFLx3_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_SDFLx3_ASAP7_75t_R%NET061 VSS N_MM29_d N_MM32_s N_NET061_1
+ PM_SDFLx3_ASAP7_75t_R%NET061
cc_1 N_NET061_1 N_MM27_g 0.0173504f
cc_2 N_NET061_1 N_MM30_g 0.0172405f
x_PM_SDFLx3_ASAP7_75t_R%noxref_33 VSS N_noxref_33_1
+ PM_SDFLx3_ASAP7_75t_R%noxref_33
cc_3 N_noxref_33_1 N_MM0_g 0.00129969f
cc_4 N_noxref_33_1 N_SEN_3 0.00192066f
cc_5 N_noxref_33_1 N_SEN_10 0.0374846f
cc_6 N_noxref_33_1 N_noxref_31_1 0.00745852f
cc_7 N_noxref_33_1 N_noxref_32_1 0.000452482f
x_PM_SDFLx3_ASAP7_75t_R%noxref_34 VSS N_noxref_34_1
+ PM_SDFLx3_ASAP7_75t_R%noxref_34
cc_8 N_noxref_34_1 N_MM0_g 0.00135268f
cc_9 N_noxref_34_1 N_SEN_3 0.000116022f
cc_10 N_noxref_34_1 N_SEN_4 0.000411435f
cc_11 N_noxref_34_1 N_SEN_11 0.0373254f
cc_12 N_noxref_34_1 N_noxref_31_1 0.000462323f
cc_13 N_noxref_34_1 N_noxref_32_1 0.00775511f
cc_14 N_noxref_34_1 N_noxref_33_1 0.00119887f
x_PM_SDFLx3_ASAP7_75t_R%noxref_35 VSS N_noxref_35_1
+ PM_SDFLx3_ASAP7_75t_R%noxref_35
cc_15 N_noxref_35_1 N_MM24@2_g 0.00148477f
cc_16 N_noxref_35_1 N_QN_14 0.0377351f
x_PM_SDFLx3_ASAP7_75t_R%noxref_31 VSS N_noxref_31_1
+ PM_SDFLx3_ASAP7_75t_R%noxref_31
cc_17 N_noxref_31_1 N_SEN_3 0.00180742f
cc_18 N_noxref_31_1 N_SS_10 0.0168947f
cc_19 N_noxref_31_1 N_MM14_g 0.00572046f
x_PM_SDFLx3_ASAP7_75t_R%noxref_32 VSS N_noxref_32_1
+ PM_SDFLx3_ASAP7_75t_R%noxref_32
cc_20 N_noxref_32_1 N_SEN_4 0.000149394f
cc_21 N_noxref_32_1 N_SEN_11 0.000897361f
cc_22 N_noxref_32_1 N_SS_11 0.0169645f
cc_23 N_noxref_32_1 N_MM14_g 0.00581205f
cc_24 N_noxref_32_1 N_noxref_31_1 0.00152625f
x_PM_SDFLx3_ASAP7_75t_R%noxref_36 VSS N_noxref_36_1
+ PM_SDFLx3_ASAP7_75t_R%noxref_36
cc_25 N_noxref_36_1 N_MM24@2_g 0.00148536f
cc_26 N_noxref_36_1 N_QN_16 0.0378228f
cc_27 N_noxref_36_1 N_noxref_35_1 0.00177583f
x_PM_SDFLx3_ASAP7_75t_R%QN VSS QN N_MM24_d N_MM24@3_d N_MM24@2_d N_MM25_d
+ N_MM25@3_d N_MM25@2_d N_QN_13 N_QN_19 N_QN_3 N_QN_15 N_QN_4 N_QN_18 N_QN_1
+ N_QN_2 N_QN_16 N_QN_14 PM_SDFLx3_ASAP7_75t_R%QN
cc_28 N_QN_13 N_SH_22 0.00113276f
cc_29 N_QN_13 N_SH_2 0.000427363f
cc_30 N_QN_13 N_MM24@2_g 0.00093274f
cc_31 N_QN_13 N_SH_27 0.00060768f
cc_32 N_QN_19 N_SH_2 0.000812406f
cc_33 N_QN_3 N_MM24@2_g 0.000856681f
cc_34 N_QN_15 N_MM24_g 0.0309691f
cc_35 N_QN_4 N_MM24@2_g 0.000912787f
cc_36 N_QN_18 N_SH_22 0.00122298f
cc_37 N_QN_1 N_MM24_g 0.0021107f
cc_38 N_QN_2 N_SH_22 0.00233502f
cc_39 N_QN_2 N_MM24_g 0.0023405f
cc_40 N_QN_16 N_MM24@2_g 0.0151252f
cc_41 N_QN_15 N_SH_2 0.00674893f
cc_42 N_QN_14 N_MM24@2_g 0.0525327f
cc_43 N_QN_13 N_MM24@3_g 0.0372853f
cc_44 N_QN_13 N_MM24_g 0.0682103f
x_PM_SDFLx3_ASAP7_75t_R%D VSS D N_MM30_g N_D_1 N_D_5 PM_SDFLx3_ASAP7_75t_R%D
cc_45 N_MM30_g N_SEN_16 0.000481842f
cc_46 N_MM30_g N_SEN_1 0.000865616f
cc_47 N_D_1 N_SEN_1 0.00120732f
cc_48 N_D_5 N_SEN_14 0.00159242f
cc_49 N_D N_SEN_12 0.0021517f
cc_50 N_MM30_g N_MM27_g 0.00504614f
x_PM_SDFLx3_ASAP7_75t_R%NET062 VSS N_MM26_d N_MM5_s N_NET062_7 N_NET062_9
+ N_NET062_1 N_NET062_11 N_NET062_12 N_NET062_10 N_NET062_8 N_NET062_2
+ PM_SDFLx3_ASAP7_75t_R%NET062
cc_51 N_NET062_7 N_SE_1 0.00126014f
cc_52 N_NET062_9 N_SE_10 0.000665467f
cc_53 N_NET062_1 N_SE_8 0.000836842f
cc_54 N_NET062_11 N_SE_7 0.0012823f
cc_55 N_NET062_12 N_SE_10 0.00135788f
cc_56 N_NET062_1 N_MM31_g 0.00159009f
cc_57 N_NET062_11 N_SE_8 0.00389037f
cc_58 N_NET062_10 N_SE_13 0.00437359f
cc_59 N_NET062_7 N_MM31_g 0.034181f
cc_60 N_NET062_10 N_SEN_12 0.000325622f
cc_61 N_NET062_10 N_SEN_16 0.000381283f
cc_62 N_NET062_11 N_SEN_12 0.00109722f
cc_63 N_NET062_10 N_SEN_14 0.00547736f
cc_64 N_NET062_8 N_SI_1 0.00130049f
cc_65 N_NET062_2 N_MM3_g 0.00153465f
cc_66 N_NET062_8 N_MM3_g 0.0349087f
x_PM_SDFLx3_ASAP7_75t_R%noxref_29 VSS N_noxref_29_1
+ PM_SDFLx3_ASAP7_75t_R%noxref_29
cc_67 N_noxref_29_1 N_MM31_g 0.00147391f
cc_68 N_noxref_29_1 N_CLKB_14 0.000676707f
cc_69 N_noxref_29_1 N_PU1_8 0.0360702f
cc_70 N_noxref_29_1 N_noxref_26_1 0.000466525f
cc_71 N_noxref_29_1 N_noxref_27_1 0.00771767f
cc_72 N_noxref_29_1 N_noxref_28_1 0.00123961f
x_PM_SDFLx3_ASAP7_75t_R%noxref_28 VSS N_noxref_28_1
+ PM_SDFLx3_ASAP7_75t_R%noxref_28
cc_73 N_noxref_28_1 N_MM31_g 0.00165253f
cc_74 N_noxref_28_1 N_CLKB_13 0.000612844f
cc_75 N_noxref_28_1 N_NET062_7 0.0360283f
cc_76 N_noxref_28_1 N_noxref_26_1 0.00769512f
cc_77 N_noxref_28_1 N_noxref_27_1 0.000469727f
x_PM_SDFLx3_ASAP7_75t_R%SE VSS SE N_MM31_g N_MM0_g N_SE_9 N_SE_13 N_SE_8
+ N_SE_12 N_SE_1 N_SE_2 N_SE_10 N_SE_7 N_SE_11 PM_SDFLx3_ASAP7_75t_R%SE
x_PM_SDFLx3_ASAP7_75t_R%CLK VSS CLK N_MM20_g N_CLK_4 N_CLK_6 N_CLK_1 N_CLK_5
+ PM_SDFLx3_ASAP7_75t_R%CLK
x_PM_SDFLx3_ASAP7_75t_R%NET063 VSS N_MM31_s N_MM27_d N_MM30_d N_MM3_s
+ N_NET063_9 N_NET063_7 N_NET063_1 N_NET063_2 N_NET063_8
+ PM_SDFLx3_ASAP7_75t_R%NET063
cc_78 N_NET063_9 N_CLKN_35 0.00296013f
cc_79 N_NET063_7 N_SE_1 0.000976129f
cc_80 N_NET063_9 N_SE_8 0.000729058f
cc_81 N_NET063_1 N_MM31_g 0.000834141f
cc_82 N_NET063_7 N_MM31_g 0.0328594f
cc_83 N_NET063_7 N_SEN_1 0.000919033f
cc_84 N_NET063_1 N_MM27_g 0.000850859f
cc_85 N_NET063_9 N_SEN_12 0.00208069f
cc_86 N_NET063_7 N_MM27_g 0.0329447f
cc_87 N_NET063_2 N_MM30_g 0.00086414f
cc_88 N_NET063_9 N_D 0.00224335f
cc_89 N_NET063_8 N_MM30_g 0.0339626f
cc_90 N_NET063_9 N_SI_4 0.00061549f
cc_91 N_NET063_8 N_SI_1 0.000776146f
cc_92 N_NET063_2 N_MM3_g 0.000815023f
cc_93 N_NET063_8 N_MM3_g 0.0335002f
cc_94 N_NET063_2 N_PU1_11 0.000546842f
cc_95 N_NET063_7 N_PU1_8 0.00110342f
cc_96 N_NET063_8 N_PU1_9 0.000553893f
cc_97 N_NET063_1 N_PU1_11 0.000596544f
cc_98 N_NET063_8 N_PU1_2 0.00129778f
cc_99 N_NET063_2 N_PU1_2 0.00160893f
cc_100 N_NET063_1 N_PU1_1 0.00302503f
cc_101 N_NET063_9 N_PU1_11 0.0128284f
x_PM_SDFLx3_ASAP7_75t_R%SEN VSS N_MM27_g N_MM0_d N_MM2_d N_SEN_3 N_SEN_4
+ N_SEN_13 N_SEN_14 N_SEN_1 N_SEN_15 N_SEN_11 N_SEN_10 N_SEN_12 N_SEN_16
+ PM_SDFLx3_ASAP7_75t_R%SEN
cc_102 N_SEN_3 N_SE_9 0.000160442f
cc_103 N_SEN_4 N_SE_9 0.000167851f
cc_104 N_SEN_13 N_SE_9 0.00807423f
cc_105 N_SEN_14 N_SE_13 0.000247294f
cc_106 N_SEN_1 N_SE_8 0.000309112f
cc_107 N_SEN_13 N_SE_12 0.000345458f
cc_108 N_SEN_15 N_SE_9 0.000409821f
cc_109 N_SEN_11 N_MM0_g 0.0159389f
cc_110 N_SEN_10 N_MM0_g 0.05362f
cc_111 N_SEN_1 N_SE_1 0.00125681f
cc_112 N_SEN_12 N_SE_13 0.000479967f
cc_113 N_SEN_13 N_SE_13 0.000508708f
cc_114 N_SEN_4 N_SE_2 0.000687367f
cc_115 N_SEN_4 N_MM0_g 0.0013466f
cc_116 N_SEN_12 N_SE_8 0.00168423f
cc_117 N_SEN_3 N_MM0_g 0.00173632f
cc_118 N_SEN_11 N_SE_2 0.00177179f
cc_119 N_MM27_g N_MM31_g 0.00330887f
cc_120 N_SEN_16 N_SE_13 0.0666113f
x_PM_SDFLx3_ASAP7_75t_R%PD2 VSS N_MM10_s N_MM11_d N_PD2_4 N_PD2_5 N_PD2_1
+ PM_SDFLx3_ASAP7_75t_R%PD2
cc_121 N_PD2_4 N_CLKN_29 8.52576e-20
cc_122 N_PD2_4 N_CLKN_10 0.000126144f
cc_123 N_PD2_4 N_CLKN_3 0.000277545f
cc_124 N_PD2_5 N_CLKN_10 0.00167232f
cc_125 N_PD2_1 N_MM9_g 0.00209534f
cc_126 N_PD2_5 N_MM9_g 0.00734593f
cc_127 N_PD2_4 N_MM9_g 0.0237369f
cc_128 N_PD2_4 N_MM10_g 0.0150074f
cc_129 N_PD2_5 N_MM11_g 0.0148527f
cc_130 N_PD2_4 N_MH_14 0.000321573f
cc_131 N_PD2_4 N_MH_3 0.000612684f
cc_132 N_PD2_1 N_MH_14 0.0034933f
x_PM_SDFLx3_ASAP7_75t_R%PD3 VSS N_MM9_s N_MM8_d N_PD3_1
+ PM_SDFLx3_ASAP7_75t_R%PD3
cc_133 N_PD3_1 N_MM9_g 0.00777391f
cc_134 N_PD3_1 N_MM11_g 0.0078334f
x_PM_SDFLx3_ASAP7_75t_R%PD5 VSS N_MM17_s N_MM16_d N_PD5_1 N_PD5_5 N_PD5_4
+ PM_SDFLx3_ASAP7_75t_R%PD5
cc_135 N_PD5_1 N_MM18_g 0.000757693f
cc_136 N_PD5_5 N_MM18_g 0.00693413f
cc_137 N_PD5_4 N_MM18_g 0.0239667f
cc_138 N_PD5_4 N_MM17_g 0.0152567f
cc_139 N_PD5_1 N_MM16_g 0.00089213f
cc_140 N_PD5_5 N_MM16_g 0.0155961f
cc_141 N_PD5_1 N_SH_15 0.000514941f
cc_142 N_PD5_1 N_SH_17 0.000490506f
cc_143 N_PD5_1 N_SH_18 0.000570964f
cc_144 N_PD5_4 N_SH_5 0.000658152f
cc_145 N_PD5_1 N_SH_24 0.00238086f
x_PM_SDFLx3_ASAP7_75t_R%SI VSS SI N_MM3_g N_SI_5 N_SI_6 N_SI_7 N_SI_1 N_SI_4
+ PM_SDFLx3_ASAP7_75t_R%SI
cc_146 N_SI_5 N_CLKN_2 0.000464688f
cc_147 N_SI_5 N_MM1_g 7.54599e-20
cc_148 N_SI_5 N_CLKN_35 0.00103845f
cc_149 N_SI_6 N_CLKN_35 0.000321601f
cc_150 N_SI_7 N_CLKN_28 0.000820405f
cc_151 N_SI_6 N_CLKN_34 0.000920438f
cc_152 N_SI_5 N_CLKN_28 0.00259564f
cc_153 N_SI_1 N_MM30_g 0.000900113f
cc_154 N_SI_4 N_D_5 0.00100819f
cc_155 N_MM3_g N_MM30_g 0.00404453f
x_PM_SDFLx3_ASAP7_75t_R%PD4 VSS N_MM18_s N_MM19_d N_PD4_1
+ PM_SDFLx3_ASAP7_75t_R%PD4
cc_156 N_PD4_1 N_MM18_g 0.00783214f
cc_157 N_PD4_1 N_MM16_g 0.00773625f
x_PM_SDFLx3_ASAP7_75t_R%noxref_26 VSS N_noxref_26_1
+ PM_SDFLx3_ASAP7_75t_R%noxref_26
cc_158 N_noxref_26_1 N_CLKN_1 0.000129154f
cc_159 N_noxref_26_1 N_MM22_g 0.00339694f
cc_160 N_noxref_26_1 N_CLKB_5 0.000434421f
cc_161 N_noxref_26_1 N_CLKB_13 0.0271823f
cc_162 N_noxref_26_1 N_NET062_7 0.000552964f
x_PM_SDFLx3_ASAP7_75t_R%PU1 VSS N_MM31_d N_MM3_d N_MM1_s N_PU1_10 N_PU1_2
+ N_PU1_11 N_PU1_8 N_PU1_1 N_PU1_9 PM_SDFLx3_ASAP7_75t_R%PU1
cc_163 N_PU1_10 N_CLKN_28 0.000382004f
cc_164 N_PU1_10 N_MM22_g 3.38254e-20
cc_165 N_PU1_10 N_CLKN_35 8.76681e-20
cc_166 N_PU1_10 N_CLKN_2 0.00101404f
cc_167 N_PU1_10 N_CLKN_34 0.000340781f
cc_168 N_PU1_2 N_MM1_g 0.00159172f
cc_169 N_PU1_11 N_CLKN_35 0.00339974f
cc_170 N_PU1_10 N_MM1_g 0.0339454f
cc_171 N_PU1_8 N_SE_8 0.000751958f
cc_172 N_PU1_8 N_SE_1 0.0010048f
cc_173 N_PU1_1 N_MM31_g 0.00131636f
cc_174 N_PU1_8 N_MM31_g 0.0341575f
cc_175 N_PU1_2 N_SI_5 0.000639659f
cc_176 N_PU1_9 N_SI_1 0.00143753f
cc_177 N_PU1_2 N_SI_6 0.00293894f
cc_178 N_PU1_11 N_SI_6 0.00314952f
cc_179 N_PU1_9 N_MM3_g 0.0350635f
cc_180 N_PU1_2 N_MH_3 0.00118998f
cc_181 N_PU1_2 N_MH_12 0.00291013f
x_PM_SDFLx3_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_SDFLx3_ASAP7_75t_R%noxref_24
cc_182 N_noxref_24_1 N_MM20_g 0.00368531f
cc_183 N_noxref_24_1 N_CLKN_31 3.2883e-20
cc_184 N_noxref_24_1 N_CLKN_8 0.000549624f
cc_185 N_noxref_24_1 N_CLKN_9 4.41927e-20
cc_186 N_noxref_24_1 N_CLKN_30 5.4907e-20
cc_187 N_noxref_24_1 N_CLKN_23 0.000386523f
cc_188 N_noxref_24_1 N_CLKN_21 0.0275622f
x_PM_SDFLx3_ASAP7_75t_R%noxref_27 VSS N_noxref_27_1
+ PM_SDFLx3_ASAP7_75t_R%noxref_27
cc_189 N_noxref_27_1 N_CLKN_1 0.000129336f
cc_190 N_noxref_27_1 N_MM22_g 0.00342806f
cc_191 N_noxref_27_1 N_CLKB_6 0.000367361f
cc_192 N_noxref_27_1 N_CLKB_14 0.0271354f
cc_193 N_noxref_27_1 N_PU1_8 0.000589532f
cc_194 N_noxref_27_1 N_noxref_26_1 0.00148611f
x_PM_SDFLx3_ASAP7_75t_R%SS VSS N_MM16_g N_MM14_d N_MM15_d N_SS_13 N_SS_15
+ N_SS_14 N_SS_17 N_SS_16 N_SS_12 N_SS_3 N_SS_4 N_SS_1 N_SS_10 N_SS_11
+ PM_SDFLx3_ASAP7_75t_R%SS
cc_195 N_MM16_g N_CLKN_10 0.00067785f
cc_196 N_MM16_g N_CLKN_5 0.000426619f
cc_197 N_MM16_g N_MM18_g 0.0133637f
cc_198 N_SS_13 N_SE_13 0.000905372f
cc_199 N_SS_15 N_SE_13 0.00322852f
cc_200 N_SS_14 N_SEN_3 0.0015797f
cc_201 N_SS_14 N_SEN_11 0.000119235f
cc_202 N_SS_14 N_SEN_15 0.000121753f
cc_203 N_SS_14 N_SEN_4 0.00026012f
cc_204 N_SS_13 N_SEN_16 0.000361395f
cc_205 N_SS_17 N_SEN_13 0.000429155f
cc_206 N_SS_16 N_SEN_15 0.000775661f
cc_207 N_SS_12 N_SEN_16 0.00262143f
cc_208 N_SS_14 N_SEN_13 0.00877126f
x_PM_SDFLx3_ASAP7_75t_R%MS VSS N_MM11_g N_MM6_d N_MM12_d N_MM7_d N_MM13_d
+ N_MS_3 N_MS_15 N_MS_13 N_MS_12 N_MS_1 N_MS_17 N_MS_11 N_MS_4 N_MS_18 N_MS_19
+ N_MS_14 N_MS_16 PM_SDFLx3_ASAP7_75t_R%MS
cc_209 N_MS_3 N_CLKN_29 0.00014273f
cc_210 N_MS_3 N_CLKN_10 0.000652432f
cc_211 N_MS_3 N_CLKN_3 9.25654e-20
cc_212 N_MS_3 N_CLKN_35 0.000141525f
cc_213 N_MS_15 N_CLKN_29 0.000281055f
cc_214 N_MS_13 N_MM12_g 0.00786932f
cc_215 N_MS_15 N_CLKN_10 0.000361999f
cc_216 N_MS_12 N_MM12_g 0.00781547f
cc_217 N_MS_1 N_MM9_g 0.000704144f
cc_218 N_MS_17 N_CLKN_10 0.00154171f
cc_219 N_MS_11 N_MM12_g 0.006509f
cc_220 N_MS_4 N_MM12_g 0.00257216f
cc_221 N_MS_4 N_CLKN_10 0.00639206f
cc_222 N_MM11_g N_MM9_g 0.0141709f
cc_223 N_MS_3 N_MM12_g 0.0259821f
cc_224 N_MS_18 N_SEN_16 0.00092209f
cc_225 N_MS_19 N_SEN_16 0.00303751f
cc_226 N_MS_13 N_MM10_g 0.000137844f
cc_227 N_MS_13 N_CLKB_22 0.000349468f
cc_228 N_MS_13 N_CLKB_18 0.000180975f
cc_229 N_MS_13 N_CLKB_2 0.000222252f
cc_230 N_MS_17 N_CLKB_18 0.0045503f
cc_231 N_MS_17 N_CLKB_2 0.000289706f
cc_232 N_MS_19 N_CLKB_18 0.000418989f
cc_233 N_MS_18 N_CLKB_22 0.00167154f
cc_234 N_MS_13 N_MM17_g 0.0155691f
x_PM_SDFLx3_ASAP7_75t_R%PD1 VSS N_MM32_d N_MM5_d N_MM4_s N_PD1_8 N_PD1_2
+ N_PD1_9 N_PD1_7 N_PD1_1 PM_SDFLx3_ASAP7_75t_R%PD1
cc_235 N_PD1_8 N_CLKN_28 0.000153144f
cc_236 N_PD1_8 N_CLKN_2 0.00111457f
cc_237 N_PD1_2 N_MM1_g 0.00116675f
cc_238 N_PD1_9 N_CLKN_28 0.0023646f
cc_239 N_PD1_8 N_MM1_g 0.0355837f
cc_240 N_PD1_9 N_SE_13 0.00227176f
cc_241 N_PD1_9 N_MM27_g 0.000310043f
cc_242 N_PD1_9 N_SEN_12 0.000106326f
cc_243 N_PD1_9 N_SEN_14 0.000544255f
cc_244 N_PD1_9 N_SEN_16 0.00389303f
cc_245 N_PD1_7 N_D_1 0.000881032f
cc_246 N_PD1_1 N_MM30_g 0.00126293f
cc_247 N_PD1_9 N_D_5 0.00271986f
cc_248 N_PD1_7 N_MM30_g 0.034257f
cc_249 N_PD1_9 N_SI_4 0.000432312f
cc_250 N_PD1_1 N_MM3_g 0.000757368f
cc_251 N_PD1_7 N_SI_1 0.000820498f
cc_252 N_PD1_9 N_SI_7 0.00251194f
cc_253 N_PD1_7 N_MM3_g 0.0334678f
cc_254 N_PD1_8 N_CLKB_1 0.000897693f
cc_255 N_PD1_9 N_CLKB_17 0.000742715f
cc_256 N_PD1_2 N_MM10_g 0.000866334f
cc_257 N_PD1_9 N_CLKB_22 0.000909773f
cc_258 N_PD1_8 N_MM10_g 0.0327428f
cc_259 N_PD1_8 N_MH_10 0.00114799f
cc_260 N_PD1_9 N_MH_15 0.000948676f
cc_261 N_PD1_2 N_MH_4 0.00367732f
cc_262 N_PD1_7 N_NET062_10 0.000583347f
cc_263 N_PD1_9 N_NET062_2 0.000634346f
cc_264 N_PD1_7 N_NET062_8 0.000642412f
cc_265 N_PD1_1 N_NET062_2 0.00381327f
cc_266 N_PD1_9 N_NET062_10 0.00907347f
x_PM_SDFLx3_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_SDFLx3_ASAP7_75t_R%noxref_25
cc_267 N_noxref_25_1 N_MM20_g 0.00368231f
cc_268 N_noxref_25_1 N_CLKN_9 0.00053883f
cc_269 N_noxref_25_1 N_CLKN_8 4.38889e-20
cc_270 N_noxref_25_1 N_CLKN_32 5.43516e-20
cc_271 N_noxref_25_1 N_CLKN_24 7.69572e-20
cc_272 N_noxref_25_1 N_CLKN_31 9.32278e-20
cc_273 N_noxref_25_1 N_CLKN_23 0.000273893f
cc_274 N_noxref_25_1 N_CLKN_22 0.0275164f
cc_275 N_noxref_25_1 N_noxref_24_1 0.00204652f
x_PM_SDFLx3_ASAP7_75t_R%noxref_30 VSS N_noxref_30_1
+ PM_SDFLx3_ASAP7_75t_R%noxref_30
cc_276 N_noxref_30_1 N_CLKN_2 0.000184852f
cc_277 N_noxref_30_1 N_MM1_g 0.0107985f
cc_278 N_noxref_30_1 N_MM3_g 0.00149574f
cc_279 N_noxref_30_1 N_SI_1 0.00244743f
cc_280 N_noxref_30_1 N_PU1_2 0.00115938f
cc_281 N_noxref_30_1 N_PU1_10 0.0161887f
cc_282 N_noxref_30_1 N_PU1_9 0.0553152f
cc_283 N_noxref_30_1 N_NET062_8 0.0371383f
x_PM_SDFLx3_ASAP7_75t_R%MH VSS N_MM7_g N_MM4_d N_MM9_d N_MM1_d N_MM10_d N_MH_10
+ N_MH_3 N_MH_21 N_MH_17 N_MH_1 N_MH_4 N_MH_12 N_MH_14 N_MH_18 N_MH_20 N_MH_16
+ N_MH_19 N_MH_15 PM_SDFLx3_ASAP7_75t_R%MH
cc_284 N_MH_10 N_CLKN_28 0.000122535f
cc_285 N_MH_10 N_CLKN_29 0.000340718f
cc_286 N_MH_10 N_MM1_g 0.000427921f
cc_287 N_MH_10 N_CLKN_2 0.000202834f
cc_288 N_MH_3 N_CLKN_28 0.000340051f
cc_289 N_MH_3 N_CLKN_34 0.00035907f
cc_290 N_MH_21 N_CLKN_29 0.000403666f
cc_291 N_MH_17 N_CLKN_29 0.00607769f
cc_292 N_MH_17 N_CLKN_3 0.000496978f
cc_293 N_MH_1 N_CLKN_10 0.00208349f
cc_294 N_MH_4 N_MM9_g 0.000633049f
cc_295 N_MH_12 N_CLKN_2 0.000667055f
cc_296 N_MH_17 N_CLKN_10 0.000773147f
cc_297 N_MH_14 N_CLKN_35 0.00140651f
cc_298 N_MH_18 N_CLKN_29 0.00149849f
cc_299 N_MH_3 N_MM1_g 0.00156193f
cc_300 N_MH_14 N_CLKN_34 0.00371753f
cc_301 N_MM7_g N_CLKN_10 0.00508109f
cc_302 N_MH_12 N_MM1_g 0.0329691f
cc_303 N_MM7_g N_MM12_g 0.0127256f
cc_304 N_MH_10 N_MM9_g 0.0361318f
cc_305 N_MH_10 N_CLKB_17 0.000251771f
cc_306 N_MH_10 N_CLKB_2 0.000109666f
cc_307 N_MH_10 N_MM17_g 0.000136877f
cc_308 N_MH_10 N_CLKB_21 0.000293637f
cc_309 N_MH_20 N_CLKB_21 0.000318499f
cc_310 N_MH_14 N_CLKB_21 0.000451281f
cc_311 N_MH_12 N_MM10_g 0.0163537f
cc_312 N_MH_16 N_CLKB_17 0.000526618f
cc_313 N_MH_3 N_CLKB_1 0.000604473f
cc_314 N_MH_4 N_CLKB_17 0.000807397f
cc_315 N_MH_4 N_MM10_g 0.00111016f
cc_316 N_MH_3 N_MM10_g 0.00122353f
cc_317 N_MH_10 N_CLKB_1 0.00160692f
cc_318 N_MH_17 N_CLKB_21 0.00205839f
cc_319 N_MH_18 N_CLKB_22 0.00250251f
cc_320 N_MH_10 N_MM10_g 0.0526533f
cc_321 N_MH_19 N_MS_18 0.000266998f
cc_322 N_MH_4 N_MS_1 0.000360052f
cc_323 N_MH_18 N_MS_19 0.000373564f
cc_324 N_MH_18 N_MS_1 0.000662176f
cc_325 N_MM7_g N_MS_3 0.000936785f
cc_326 N_MH_18 N_MS_17 0.000996322f
cc_327 N_MH_1 N_MS_14 0.00100229f
cc_328 N_MH_1 N_MS_1 0.00130115f
cc_329 N_MM7_g N_MS_12 0.00631888f
cc_330 N_MM7_g N_MS_1 0.0024104f
cc_331 N_MM7_g N_MS_11 0.00638861f
cc_332 N_MH_18 N_MS_14 0.0045882f
cc_333 N_MH_16 N_MS_18 0.00496962f
cc_334 N_MM7_g N_MM11_g 0.0293331f
x_PM_SDFLx3_ASAP7_75t_R%CLKB VSS N_MM10_g N_MM17_g N_MM23_d N_MM22_d N_CLKB_13
+ N_CLKB_22 N_CLKB_16 N_CLKB_5 N_CLKB_19 N_CLKB_15 N_CLKB_6 N_CLKB_20 N_CLKB_14
+ N_CLKB_17 N_CLKB_18 N_CLKB_2 N_CLKB_1 N_CLKB_21 PM_SDFLx3_ASAP7_75t_R%CLKB
cc_335 N_CLKB_13 N_CLK_5 7.99986e-20
cc_336 N_CLKB_22 N_CLK_5 0.000120717f
cc_337 N_CLKB_16 N_CLK_5 0.000545781f
cc_338 N_CLKB_5 N_CLK_5 0.000386667f
cc_339 N_CLKB_19 N_CLK_5 0.00220898f
cc_340 N_CLKB_22 N_CLKN_10 2.85014e-20
cc_341 N_CLKB_22 N_CLKN_8 3.26977e-20
cc_342 N_CLKB_22 N_CLKN_25 3.59144e-20
cc_343 N_CLKB_22 N_MM22_g 4.9972e-20
cc_344 N_CLKB_5 N_CLKN_23 7.92643e-20
cc_345 N_CLKB_15 N_CLKN_26 0.00010366f
cc_346 N_CLKB_19 N_CLKN_27 0.000123067f
cc_347 N_CLKB_6 N_CLKN_33 0.000176973f
cc_348 N_MM17_g N_CLKN_5 0.000208159f
cc_349 N_CLKB_20 N_CLKN_33 0.000230779f
cc_350 N_CLKB_22 N_CLKN_29 0.000676953f
cc_351 N_CLKB_22 N_CLKN_28 0.000327609f
cc_352 N_CLKB_15 N_CLKN_27 0.000370527f
cc_353 N_CLKB_13 N_MM22_g 0.0386446f
cc_354 N_CLKB_14 N_MM22_g 0.0111649f
cc_355 N_CLKB_17 N_CLKN_35 0.000478614f
cc_356 N_CLKB_18 N_CLKN_10 0.000531969f
cc_357 N_CLKB_16 N_CLKN_1 0.000556157f
cc_358 N_MM10_g N_CLKN_3 0.000560153f
cc_359 N_CLKB_5 N_MM22_g 0.000594332f
cc_360 N_CLKB_16 N_CLKN_35 0.000617175f
cc_361 N_CLKB_2 N_CLKN_10 0.0027913f
cc_362 N_CLKB_14 N_CLKN_1 0.000776391f
cc_363 N_CLKB_6 N_MM22_g 0.000849536f
cc_364 N_CLKB_1 N_CLKN_2 0.00222254f
cc_365 N_CLKB_21 N_CLKN_34 0.00165668f
cc_366 N_CLKB_17 N_CLKN_28 0.00265567f
cc_367 N_CLKB_15 N_CLKN_33 0.00352324f
cc_368 N_MM10_g N_MM9_g 0.00370558f
cc_369 N_CLKB_16 N_CLKN_27 0.00487527f
cc_370 N_MM17_g N_CLKN_10 0.00493103f
cc_371 N_MM17_g N_MM18_g 0.00578276f
cc_372 N_MM10_g N_MM1_g 0.00704312f
cc_373 N_MM17_g N_MM12_g 0.0182761f
cc_374 N_CLKB_22 N_CLKN_35 0.0446429f
cc_375 N_CLKB_16 N_SE_1 5.26109e-20
cc_376 N_CLKB_5 N_SE_10 5.47477e-20
cc_377 N_CLKB_5 N_SE_7 0.000170428f
cc_378 N_CLKB_16 N_SE_7 0.00331576f
cc_379 N_CLKB_18 N_SE_13 0.000499861f
cc_380 N_CLKB_19 N_SE_10 0.00196725f
cc_381 N_CLKB_22 N_SE_13 0.0023571f
cc_382 N_CLKB_22 N_SE_8 0.00357592f
cc_383 N_CLKB_16 N_SE_11 0.00678176f
cc_384 N_CLKB_17 N_SEN_16 0.000503602f
cc_385 N_CLKB_22 N_SEN_12 0.00413685f
cc_386 N_CLKB_18 N_SEN_16 0.00281087f
cc_387 N_CLKB_22 N_SEN_16 0.00995472f
cc_388 N_CLKB_22 N_SI_4 0.00248601f
x_PM_SDFLx3_ASAP7_75t_R%CLKN VSS N_MM22_g N_MM1_g N_MM9_g N_MM12_g N_MM18_g
+ N_MM20_d N_MM21_d N_CLKN_30 N_CLKN_27 N_CLKN_26 N_CLKN_31 N_CLKN_8 N_CLKN_22
+ N_CLKN_21 N_CLKN_33 N_CLKN_9 N_CLKN_1 N_CLKN_35 N_CLKN_25 N_CLKN_23 N_CLKN_2
+ N_CLKN_28 N_CLKN_34 N_CLKN_10 N_CLKN_5 N_CLKN_29 N_CLKN_3 N_CLKN_32 N_CLKN_24
+ PM_SDFLx3_ASAP7_75t_R%CLKN
cc_389 N_CLKN_30 N_MM20_g 5.92433e-20
cc_390 N_CLKN_27 N_MM20_g 7.17161e-20
cc_391 N_CLKN_26 N_MM20_g 8.98024e-20
cc_392 N_CLKN_31 N_MM20_g 9.82155e-20
cc_393 N_CLKN_8 N_MM20_g 0.00111234f
cc_394 N_CLKN_22 N_MM20_g 0.0112003f
cc_395 N_CLKN_21 N_MM20_g 0.0112112f
cc_396 N_CLKN_33 N_MM20_g 0.000355378f
cc_397 N_CLKN_31 N_CLK_4 0.000415112f
cc_398 N_CLKN_9 N_MM20_g 0.000630561f
cc_399 N_CLKN_1 N_CLK_6 0.00063244f
cc_400 N_CLKN_35 N_CLK_4 0.000645354f
cc_401 N_CLKN_25 N_CLK_6 0.000943393f
cc_402 N_CLKN_27 N_CLK_6 0.000948166f
cc_403 N_CLKN_1 N_CLK_1 0.00348994f
cc_404 N_CLKN_23 N_CLK_4 0.00164912f
cc_405 N_CLKN_25 N_CLK_5 0.00176865f
cc_406 N_CLKN_27 N_CLK_4 0.00477924f
cc_407 N_MM22_g N_MM20_g 0.0350676f
x_PM_SDFLx3_ASAP7_75t_R%SH VSS N_MM14_g N_MM24_g N_MM24@3_g N_MM24@2_g N_MM13_s
+ N_MM18_d N_MM12_s N_MM17_d N_SH_16 N_SH_17 N_SH_23 N_SH_25 N_SH_15 N_SH_6
+ N_SH_20 N_SH_18 N_SH_19 N_SH_5 N_SH_22 N_SH_24 N_SH_2 N_SH_27 N_SH_1 N_SH_21
+ N_SH_26 PM_SDFLx3_ASAP7_75t_R%SH
cc_408 N_SH_16 N_CLKN_10 8.49463e-20
cc_409 N_SH_17 N_CLKN_35 9.66047e-20
cc_410 N_SH_23 N_CLKN_10 0.000196768f
cc_411 N_SH_25 N_CLKN_10 0.000203975f
cc_412 N_SH_15 N_MM12_g 0.00680288f
cc_413 N_SH_6 N_CLKN_10 0.000276295f
cc_414 N_SH_20 N_CLKN_10 0.000396208f
cc_415 N_SH_18 N_CLKN_10 0.000448364f
cc_416 N_SH_19 N_CLKN_10 0.00060535f
cc_417 N_SH_16 N_CLKN_5 0.000673075f
cc_418 N_SH_6 N_MM18_g 0.00100239f
cc_419 N_SH_5 N_CLKN_10 0.00282638f
cc_420 N_SH_5 N_MM12_g 0.00948039f
cc_421 N_SH_16 N_MM18_g 0.0160733f
cc_422 N_SH_22 N_SE_12 0.000231716f
cc_423 N_SH_24 N_SE_13 0.000236329f
cc_424 N_SH_2 N_SE_2 0.00182381f
cc_425 N_SH_17 N_SE_13 0.00102453f
cc_426 N_SH_27 N_SE_13 0.00207588f
cc_427 N_SH_18 N_SE_13 0.00279298f
cc_428 N_MM24_g N_MM0_g 0.00331442f
cc_429 N_SH_22 N_SE_9 0.0060579f
cc_430 N_MM24_g N_SEN_10 5.87766e-20
cc_431 N_SH_1 N_SEN_3 0.000208718f
cc_432 N_MM24_g N_SEN_4 9.77652e-20
cc_433 N_SH_20 N_SEN_16 0.00010979f
cc_434 N_MM14_g N_SEN_3 0.000113039f
cc_435 N_SH_27 N_SEN_15 0.000117382f
cc_436 N_SH_27 N_SEN_13 0.00150773f
cc_437 N_SH_22 N_SEN_4 0.000190471f
cc_438 N_MM24_g N_SEN_3 0.000198416f
cc_439 N_SH_22 N_SEN_15 0.000261213f
cc_440 N_SH_21 N_SEN_16 0.000292155f
cc_441 N_SH_17 N_SEN_16 0.000374558f
cc_442 N_SH_27 N_SEN_16 0.00450899f
cc_443 N_SH_18 N_SEN_16 0.00610672f
cc_444 N_SH_6 N_MM17_g 0.000158318f
cc_445 N_SH_15 N_MM17_g 0.00676966f
cc_446 N_SH_16 N_MM17_g 0.00683991f
cc_447 N_SH_23 N_CLKB_18 0.000285306f
cc_448 N_SH_17 N_CLKB_18 0.000369687f
cc_449 N_SH_25 N_CLKB_18 0.000402567f
cc_450 N_SH_19 N_CLKB_18 0.000466758f
cc_451 N_SH_18 N_CLKB_2 0.000570191f
cc_452 N_SH_5 N_CLKB_2 0.000576027f
cc_453 N_SH_27 N_CLKB_22 0.000761171f
cc_454 N_SH_17 N_CLKB_22 0.00106654f
cc_455 N_SH_18 N_CLKB_18 0.00451947f
cc_456 N_SH_5 N_MM17_g 0.0183312f
cc_457 N_SH_19 N_MS_3 9.84549e-20
cc_458 N_SH_23 N_MS_3 0.000179155f
cc_459 N_SH_16 N_MS_3 0.000436412f
cc_460 N_SH_6 N_MS_3 0.000220896f
cc_461 N_SH_15 N_MS_3 0.000232021f
cc_462 N_SH_15 N_MS_11 0.000234022f
cc_463 N_SH_23 N_MS_4 0.000335655f
cc_464 N_SH_6 N_MS_4 0.000424812f
cc_465 N_SH_17 N_MS_16 0.00043823f
cc_466 N_SH_23 N_MS_17 0.000518386f
cc_467 N_SH_16 N_MS_4 0.00059315f
cc_468 N_SH_17 N_MS_19 0.00132439f
cc_469 N_SH_5 N_MS_3 0.00373302f
cc_470 N_SH_19 N_MM16_g 9.92275e-20
cc_471 N_SH_21 N_SS_13 0.000310651f
cc_472 N_MM14_g N_SS_3 0.000322169f
cc_473 N_MM14_g N_SS_4 0.000425437f
cc_474 N_SH_24 N_SS_15 0.000580125f
cc_475 N_SH_26 N_SS_16 0.000623015f
cc_476 N_SH_26 N_SS_14 0.000697123f
cc_477 N_SH_18 N_SS_1 0.000810777f
cc_478 N_SH_1 N_SS_14 0.000950422f
cc_479 N_MM14_g N_SS_1 0.00111309f
cc_480 N_SH_1 N_MM16_g 0.00129928f
cc_481 N_SH_20 N_SS_12 0.00154842f
cc_482 N_SH_27 N_SS_14 0.0017411f
cc_483 N_MM14_g N_SS_10 0.00649524f
cc_484 N_MM14_g N_SS_11 0.0066006f
cc_485 N_SH_18 N_SS_12 0.00462671f
cc_486 N_SH_21 N_SS_14 0.00472659f
cc_487 N_MM14_g N_MM16_g 0.0300233f
*END of SDFLx3_ASAP7_75t_R.pxi
.ENDS
** Design:	SDFLx4_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "SDFLx4_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "SDFLx4_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_SDFLx4_ASAP7_75t_R%NET066 VSS 2 3 1
c1 1 VSS 0.0010093f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4860 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0675 $X2=0.4860 $Y2=0.0675
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%NET067 VSS 2 3 1
c1 1 VSS 0.00101903f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0675 $X2=0.5940 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.0675 $X2=0.5940 $Y2=0.0675
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%noxref_31 VSS 1
c1 1 VSS 0.00552771f
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%noxref_32 VSS 1
c1 1 VSS 0.00662221f
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%noxref_30 VSS 1
c1 1 VSS 0.00538347f
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.00465783f
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.00462901f
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%PD5 VSS 2 4 1
c1 1 VSS 0.00096906f
r1 4 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.2050 $Y=0.0675 $X2=1.1925 $Y2=0.0675
r2 2 1 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.1710 $Y=0.0675 $X2=1.1755 $Y2=0.0675
r3 1 3 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.1755 $Y=0.0675 $X2=1.1925 $Y2=0.0675
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%PD3 VSS 7 9 4 5 1
c1 1 VSS 0.0103267f
c2 4 VSS 0.00189632f
c3 5 VSS 0.00320808f
r1 9 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8810 $Y=0.0675 $X2=0.8785 $Y2=0.0675
r2 5 8 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8660 $Y=0.0675 $X2=0.8785 $Y2=0.0675
r3 4 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.0675 $X2=0.8080 $Y2=0.0675
r4 7 4 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.0675 $X2=0.7955 $Y2=0.0675
r5 1 5 1e-05
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%noxref_27 VSS 1
c1 1 VSS 0.00547669f
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%noxref_26 VSS 1
c1 1 VSS 0.00542658f
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%noxref_29 VSS 1
c1 1 VSS 0.0419587f
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%PD2 VSS 5 8 3 1
c1 1 VSS 0.00513574f
c2 3 VSS 0.0033196f
r1 8 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8810 $Y=0.2025 $X2=0.8785 $Y2=0.2025
r2 1 7 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8660 $Y=0.2025 $X2=0.8785 $Y2=0.2025
r3 4 1 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8540 $Y=0.2025 $X2=0.8660 $Y2=0.2025
r4 3 4 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.2025 $X2=0.8540 $Y2=0.2025
r5 5 3 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.2025 $X2=0.8495 $Y2=0.2025
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%noxref_28 VSS 1
c1 1 VSS 0.0419602f
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%noxref_35 VSS 1
c1 1 VSS 0.00960185f
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%CLK VSS 9 3 4 5 1
c1 1 VSS 0.00634971f
c2 3 VSS 0.0815005f
c3 4 VSS 0.00383859f
c4 5 VSS 0.00282093f
r1 5 8 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0720 $X2=0.0810 $Y2=0.0920
r2 7 8 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1055 $X2=0.0810 $Y2=0.0920
r3 4 7 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1170 $X2=0.0810 $Y2=0.1055
r4 9 4 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1170
r5 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r6 9 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%PD1 VSS 11 21 24 9 7 1 8 2
c1 1 VSS 0.00608278f
c2 2 VSS 0.00530152f
c3 7 VSS 0.00363401f
c4 8 VSS 0.00260088f
c5 9 VSS 0.0235483f
r1 24 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.0675 $X2=0.6625 $Y2=0.0675
r2 22 23 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6580 $Y=0.0675 $X2=0.6625 $Y2=0.0675
r3 2 22 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6460 $Y=0.0675 $X2=0.6580 $Y2=0.0675
r4 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0675 $X2=0.6460 $Y2=0.0675
r5 21 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.0675 $X2=0.6335 $Y2=0.0675
r6 2 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.0675
+ $X2=0.6480 $Y2=0.0360
r7 17 18 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6255
+ $Y=0.0360 $X2=0.6480 $Y2=0.0360
r8 16 17 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6055
+ $Y=0.0360 $X2=0.6255 $Y2=0.0360
r9 15 16 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5785
+ $Y=0.0360 $X2=0.6055 $Y2=0.0360
r10 14 15 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.0360 $X2=0.5785 $Y2=0.0360
r11 13 14 13.6416 $w=1.3e-08 $l=5.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4815
+ $Y=0.0360 $X2=0.5400 $Y2=0.0360
r12 12 13 11.5429 $w=1.3e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4815 $Y2=0.0360
r13 9 12 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4205
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r14 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4320 $Y2=0.0360
r15 11 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r16 7 10 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4340 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r17 1 7 1e-05
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%noxref_33 VSS 1
c1 1 VSS 0.00652227f
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%D VSS 12 3 7 1 10 8 9 5 4 6
c1 1 VSS 0.0045875f
c2 3 VSS 0.0448712f
c3 4 VSS 0.00214845f
c4 5 VSS 0.00208523f
c5 6 VSS 0.00792274f
c6 7 VSS 0.0016868f
c7 8 VSS 0.001432f
c8 9 VSS 0.00379314f
c9 10 VSS 0.00144808f
r1 6 9 3.59766 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4095
+ $Y=0.2340 $X2=0.3870 $Y2=0.2340
r2 9 17 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3870
+ $Y=0.2340 $X2=0.3870 $Y2=0.2160
r3 16 17 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3870
+ $Y=0.1980 $X2=0.3870 $Y2=0.2160
r4 15 16 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3870
+ $Y=0.1765 $X2=0.3870 $Y2=0.1980
r5 4 8 5.92955 $w=1.57138e-08 $l=3.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3870 $Y=0.1405 $X2=0.3870 $Y2=0.1080
r6 4 15 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.3870
+ $Y=0.1405 $X2=0.3870 $Y2=0.1765
r7 8 14 3.59766 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3870
+ $Y=0.1080 $X2=0.4095 $Y2=0.1080
r8 5 10 3.59766 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4365
+ $Y=0.1080 $X2=0.4590 $Y2=0.1080
r9 5 14 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4365
+ $Y=0.1080 $X2=0.4095 $Y2=0.1080
r10 12 7 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1215
r11 7 10 1.49895 $w=1.95333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1215 $X2=0.4590 $Y2=0.1080
r12 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r13 12 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1350
+ $X2=0.4590 $Y2=0.1350
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%SEN VSS 9 37 39 10 17 16 11 4 1 19 3 13 15 14
c1 1 VSS 0.00389951f
c2 3 VSS 0.00773635f
c3 4 VSS 0.00803669f
c4 9 VSS 0.0815925f
c5 10 VSS 0.0052757f
c6 11 VSS 0.0053002f
c7 12 VSS 0.00048153f
c8 13 VSS 0.00429212f
c9 14 VSS 0.00202619f
c10 15 VSS 0.00299899f
c11 16 VSS 0.00757265f
c12 17 VSS 0.00563737f
c13 18 VSS 0.000260661f
c14 19 VSS 0.0006056f
r1 11 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3220 $Y2=0.2025
r2 39 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r3 10 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3220 $Y2=0.0675
r4 37 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r5 4 34 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.2340
r6 3 31 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0675
+ $X2=0.3240 $Y2=0.0360
r7 34 35 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.2340 $X2=0.3375 $Y2=0.2340
r8 17 29 10.3626 $w=1.39091e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.2340 $X2=0.3510 $Y2=0.1845
r9 17 35 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.2340 $X2=0.3375 $Y2=0.2340
r10 31 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.0360 $X2=0.3375 $Y2=0.0360
r11 16 32 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.0360 $X2=0.3375 $Y2=0.0360
r12 28 29 11.5429 $w=1.3e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1845
r13 27 28 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1125 $X2=0.3510 $Y2=0.1350
r14 13 18 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0900 $X2=0.3510 $Y2=0.0720
r15 13 27 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0900 $X2=0.3510 $Y2=0.1125
r16 12 18 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0540 $X2=0.3510 $Y2=0.0720
r17 12 16 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0540 $X2=0.3510 $Y2=0.0360
r18 18 26 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0720 $X2=0.3690 $Y2=0.0720
r19 25 26 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.3980
+ $Y=0.0720 $X2=0.3690 $Y2=0.0720
r20 24 25 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4430
+ $Y=0.0720 $X2=0.3980 $Y2=0.0720
r21 14 19 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4860 $Y=0.0720 $X2=0.5130 $Y2=0.0720
r22 14 24 10.0272 $w=1.3e-08 $l=4.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.0720 $X2=0.4430 $Y2=0.0720
r23 19 23 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0720 $X2=0.5130 $Y2=0.0900
r24 15 21 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1125 $X2=0.5130 $Y2=0.1350
r25 15 23 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1125 $X2=0.5130 $Y2=0.0900
r26 9 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r27 1 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.1350
+ $X2=0.5130 $Y2=0.1350
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%noxref_36 VSS 1
c1 1 VSS 0.00476289f
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%noxref_38 VSS 1
c1 1 VSS 0.0417984f
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%noxref_39 VSS 1
c1 1 VSS 0.0418856f
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%noxref_37 VSS 1
c1 1 VSS 0.00516025f
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%noxref_40 VSS 1
c1 1 VSS 0.0423303f
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%noxref_41 VSS 1
c1 1 VSS 0.0423153f
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%PD4 VSS 7 9 4 5 1
c1 1 VSS 0.00859232f
c2 4 VSS 0.00181994f
c3 5 VSS 0.00311373f
r1 9 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.2050 $Y=0.2025 $X2=1.2025 $Y2=0.2025
r2 5 8 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.1900 $Y=0.2025 $X2=1.2025 $Y2=0.2025
r3 4 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.1195 $Y=0.2025 $X2=1.1320 $Y2=0.2025
r4 7 4 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.1170 $Y=0.2025 $X2=1.1195 $Y2=0.2025
r5 1 5 1e-05
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%QN VSS 31 24 25 35 36 44 45 48 49 14 16 15 13 18
+ 17 2 3 4 1
c1 1 VSS 0.0104529f
c2 2 VSS 0.0104827f
c3 3 VSS 0.00996555f
c4 4 VSS 0.00991764f
c5 13 VSS 0.00445942f
c6 14 VSS 0.00439616f
c7 15 VSS 0.00446345f
c8 16 VSS 0.00440916f
c9 17 VSS 0.019105f
c10 18 VSS 0.0200449f
c11 19 VSS 0.00795447f
c12 20 VSS 0.00328544f
c13 21 VSS 0.00333904f
r1 49 47 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.5830 $Y=0.2025 $X2=1.5805 $Y2=0.2025
r2 4 47 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.5660 $Y=0.2025 $X2=1.5805 $Y2=0.2025
r3 16 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.5515 $Y=0.2025 $X2=1.5660 $Y2=0.2025
r4 48 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.5490 $Y=0.2025 $X2=1.5515 $Y2=0.2025
r5 45 43 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.4750 $Y=0.2025 $X2=1.4725 $Y2=0.2025
r6 2 43 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.4580 $Y=0.2025 $X2=1.4725 $Y2=0.2025
r7 15 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.4435 $Y=0.2025 $X2=1.4580 $Y2=0.2025
r8 44 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.4410 $Y=0.2025 $X2=1.4435 $Y2=0.2025
r9 4 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.5660 $Y=0.2025
+ $X2=1.5660 $Y2=0.2340
r10 2 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.4580 $Y=0.2025
+ $X2=1.4580 $Y2=0.2340
r11 39 40 9.32759 $w=1.3e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=1.5660
+ $Y=0.2340 $X2=1.6060 $Y2=0.2340
r12 38 39 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.5120
+ $Y=0.2340 $X2=1.5660 $Y2=0.2340
r13 37 38 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.4580
+ $Y=0.2340 $X2=1.5120 $Y2=0.2340
r14 18 37 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=1.4480
+ $Y=0.2340 $X2=1.4580 $Y2=0.2340
r15 21 32 8.52248 $w=1.49091e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.6465 $Y=0.2340 $X2=1.6465 $Y2=0.1845
r16 21 40 7.67296 $w=1.54395e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.6465 $Y=0.2340 $X2=1.6060 $Y2=0.2340
r17 36 34 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.5830 $Y=0.0675 $X2=1.5805 $Y2=0.0675
r18 3 34 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.5660 $Y=0.0675 $X2=1.5805 $Y2=0.0675
r19 14 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.5515 $Y=0.0675 $X2=1.5660 $Y2=0.0675
r20 35 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.5490 $Y=0.0675 $X2=1.5515 $Y2=0.0675
r21 31 32 9.8736 $w=1.4e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=1.6465
+ $Y=0.1350 $X2=1.6465 $Y2=0.1845
r22 19 20 8.52248 $w=1.49091e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.6465 $Y=0.0855 $X2=1.6465 $Y2=0.0360
r23 31 19 9.8736 $w=1.4e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=1.6465
+ $Y=0.1350 $X2=1.6465 $Y2=0.0855
r24 3 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.5660 $Y=0.0675
+ $X2=1.5660 $Y2=0.0360
r25 20 30 7.67296 $w=1.54395e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.6465 $Y=0.0360 $X2=1.6060 $Y2=0.0360
r26 29 30 9.32759 $w=1.3e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=1.5660
+ $Y=0.0360 $X2=1.6060 $Y2=0.0360
r27 28 29 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.5120
+ $Y=0.0360 $X2=1.5660 $Y2=0.0360
r28 27 28 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.4580
+ $Y=0.0360 $X2=1.5120 $Y2=0.0360
r29 26 27 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=1.4480
+ $Y=0.0360 $X2=1.4580 $Y2=0.0360
r30 17 26 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.4455
+ $Y=0.0360 $X2=1.4480 $Y2=0.0360
r31 1 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.4580 $Y=0.0675
+ $X2=1.4580 $Y2=0.0360
r32 25 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.4750 $Y=0.0675 $X2=1.4725 $Y2=0.0675
r33 1 23 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.4580 $Y=0.0675 $X2=1.4725 $Y2=0.0675
r34 13 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.4435 $Y=0.0675 $X2=1.4580 $Y2=0.0675
r35 24 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.4410 $Y=0.0675 $X2=1.4435 $Y2=0.0675
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%SS VSS 9 28 32 1 12 10 11 3 14 4 17 16 13 15
c1 1 VSS 0.00417681f
c2 3 VSS 0.00854531f
c3 4 VSS 0.00636581f
c4 9 VSS 0.0814212f
c5 10 VSS 0.00419973f
c6 11 VSS 0.00459679f
c7 12 VSS 0.00146988f
c8 13 VSS 0.00190258f
c9 14 VSS 0.00106437f
c10 15 VSS 0.000441271f
c11 16 VSS 0.00068339f
c12 17 VSS 0.000441843f
r1 10 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.2815 $Y=0.0675 $X2=1.2940 $Y2=0.0675
r2 32 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.2790 $Y=0.0675 $X2=1.2815 $Y2=0.0675
r3 3 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.3055 $Y=0.0675
+ $X2=1.2960 $Y2=0.0900
r4 29 30 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.2960
+ $Y=0.0900 $X2=1.3095 $Y2=0.0900
r5 16 26 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.0900 $X2=1.3230 $Y2=0.1125
r6 16 30 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3230 $Y=0.0900 $X2=1.3095 $Y2=0.0900
r7 11 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.2815 $Y=0.2025 $X2=1.2940 $Y2=0.2025
r8 28 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.2790 $Y=0.2025 $X2=1.2815 $Y2=0.2025
r9 25 26 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.1350 $X2=1.3230 $Y2=0.1125
r10 14 17 4.8802 $w=1.615e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.1630 $X2=1.3230 $Y2=0.1910
r11 14 25 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.1630 $X2=1.3230 $Y2=0.1350
r12 4 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.2960 $Y=0.2025
+ $X2=1.2960 $Y2=0.1910
r13 17 24 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3230 $Y=0.1910 $X2=1.3095 $Y2=0.1910
r14 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.2960
+ $Y=0.1910 $X2=1.3095 $Y2=0.1910
r15 22 23 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.2850
+ $Y=0.1910 $X2=1.2960 $Y2=0.1910
r16 21 22 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.2625
+ $Y=0.1910 $X2=1.2850 $Y2=0.1910
r17 13 15 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.2330
+ $Y=0.1910 $X2=1.2150 $Y2=0.1910
r18 13 21 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=1.2330
+ $Y=0.1910 $X2=1.2625 $Y2=0.1910
r19 15 20 4.8802 $w=1.615e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.2150
+ $Y=0.1910 $X2=1.2150 $Y2=0.1630
r20 12 20 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.2150
+ $Y=0.1350 $X2=1.2150 $Y2=0.1630
r21 9 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=1.2150
+ $Y=0.1350 $X2=1.2150 $Y2=0.1350
r22 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.2150 $Y=0.1350
+ $X2=1.2150 $Y2=0.1350
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%MS VSS 11 35 39 41 43 13 17 4 16 15 1 5 3 12 14
c1 1 VSS 0.00368282f
c2 3 VSS 0.000124003f
c3 4 VSS 0.016431f
c4 5 VSS 0.0101133f
c5 11 VSS 0.0793699f
c6 12 VSS 0.00383245f
c7 13 VSS 0.00262836f
c8 14 VSS 0.00380846f
c9 15 VSS 0.00260116f
c10 16 VSS 0.00128675f
c11 17 VSS 0.00387603f
c12 18 VSS 0.00126737f
r1 43 42 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0430 $Y=0.2025 $X2=1.0405 $Y2=0.2025
r2 15 42 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0280 $Y=0.2025 $X2=1.0405 $Y2=0.2025
r3 14 5 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9575 $Y=0.2025 $X2=0.9700 $Y2=0.2025
r4 41 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9550 $Y=0.2025 $X2=0.9575 $Y2=0.2025
r5 5 37 5.26888 $w=6.87567e-08 $l=4.85026e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9990 $Y=0.2025 $X2=0.9985 $Y2=0.1540
r6 39 38 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.0970 $Y=0.0675 $X2=1.0945 $Y2=0.0675
r7 13 38 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.0820 $Y=0.0675 $X2=1.0945 $Y2=0.0675
r8 36 37 3.71245 $w=4.12e-08 $l=1.9e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9985 $Y=0.1350 $X2=0.9985 $Y2=0.1540
r9 3 28 3.08411 $w=6.89849e-08 $l=4.86647e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9985 $Y=0.1160 $X2=1.0025 $Y2=0.0675
r10 3 36 3.71245 $w=4.12e-08 $l=1.9e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9985 $Y=0.1160 $X2=0.9985 $Y2=0.1350
r11 12 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9575 $Y=0.0675 $X2=0.9700 $Y2=0.0675
r12 35 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9550 $Y=0.0675 $X2=0.9575 $Y2=0.0675
r13 32 13 1.22083 $w=7.72e-08 $l=1.4e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.0660 $Y=0.0675 $X2=1.0800 $Y2=0.0675
r14 31 32 1.13362 $w=7.72e-08 $l=1.3e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.0530 $Y=0.0675 $X2=1.0660 $Y2=0.0675
r15 30 31 1.13362 $w=7.72e-08 $l=1.3e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.0400 $Y=0.0675 $X2=1.0530 $Y2=0.0675
r16 29 30 0.915619 $w=7.72e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.0295 $Y=0.0675 $X2=1.0400 $Y2=0.0675
r17 28 29 2.26219 $w=7.98037e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.0025 $Y=0.0675 $X2=1.0295 $Y2=0.0675
r18 27 28 1.84983 $w=8.1e-08 $l=2.25e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9800 $Y=0.0675 $X2=1.0025 $Y2=0.0675
r19 4 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.9680 $Y=0.0675
+ $X2=0.9720 $Y2=0.0720
r20 4 27 1.02647 $w=7.84667e-08 $l=1.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9680 $Y=0.0675 $X2=0.9800 $Y2=0.0675
r21 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.9585
+ $Y=0.0720 $X2=0.9720 $Y2=0.0720
r22 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.0720 $X2=0.9585 $Y2=0.0720
r23 17 18 4.75866 $w=1.41702e-08 $l=2.72259e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9180 $Y=0.0720 $X2=0.8910 $Y2=0.0755
r24 17 24 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.0720 $X2=0.9450 $Y2=0.0720
r25 18 22 3.47612 $w=1.45278e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8910 $Y=0.0755 $X2=0.8910 $Y2=0.0935
r26 16 20 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1160 $X2=0.8910 $Y2=0.1350
r27 16 22 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1160 $X2=0.8910 $Y2=0.0935
r28 11 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.8910
+ $Y=0.1350 $X2=0.8910 $Y2=0.1350
r29 1 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8910 $Y=0.1350
+ $X2=0.8910 $Y2=0.1350
r30 5 15 1e-05
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%SH VSS 11 12 13 14 15 49 52 95 98 16 6 18 17 5 19
+ 26 20 2 24 1 28 23 21 22 27 29
c1 1 VSS 0.00593098f
c2 2 VSS 0.0203055f
c3 5 VSS 0.00719829f
c4 6 VSS 0.00789178f
c5 11 VSS 0.0812412f
c6 12 VSS 0.0821605f
c7 13 VSS 0.0813808f
c8 14 VSS 0.0812985f
c9 15 VSS 0.0821209f
c10 16 VSS 0.00619533f
c11 17 VSS 0.00583485f
c12 18 VSS 0.0298683f
c13 19 VSS 0.0143857f
c14 20 VSS 0.00343279f
c15 21 VSS 0.0110869f
c16 22 VSS 0.00429668f
c17 23 VSS 0.00425788f
c18 24 VSS 0.00321614f
c19 25 VSS 0.00358981f
c20 26 VSS 0.00167755f
c21 27 VSS 0.00505315f
c22 28 VSS 0.00146157f
c23 29 VSS 0.00478375f
r1 98 97 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0970 $Y=0.2025 $X2=1.0945 $Y2=0.2025
r2 5 97 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0820 $Y=0.2025 $X2=1.0945 $Y2=0.2025
r3 94 5 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0700 $Y=0.2025 $X2=1.0820 $Y2=0.2025
r4 17 94 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0655 $Y=0.2025 $X2=1.0700 $Y2=0.2025
r5 95 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0630 $Y=0.2025 $X2=1.0655 $Y2=0.2025
r6 5 87 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0800 $Y=0.2025
+ $X2=1.0800 $Y2=0.2340
r7 15 79 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=1.5930
+ $Y=0.1350 $X2=1.5930 $Y2=0.1350
r8 14 73 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=1.5390
+ $Y=0.1350 $X2=1.5390 $Y2=0.1350
r9 13 67 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=1.4850
+ $Y=0.1350 $X2=1.4850 $Y2=0.1350
r10 12 59 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=1.4310 $Y=0.1350 $X2=1.4310 $Y2=0.1350
r11 87 88 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.0800
+ $Y=0.2340 $X2=1.0935 $Y2=0.2340
r12 85 88 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.2340 $X2=1.0935 $Y2=0.2340
r13 84 85 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.1340
+ $Y=0.2340 $X2=1.1070 $Y2=0.2340
r14 83 84 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.2340 $X2=1.1340 $Y2=0.2340
r15 82 83 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.1880
+ $Y=0.2340 $X2=1.1610 $Y2=0.2340
r16 81 82 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.2690
+ $Y=0.2340 $X2=1.1880 $Y2=0.2340
r17 18 29 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3500 $Y=0.2340 $X2=1.3770 $Y2=0.2340
r18 18 81 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.3500
+ $Y=0.2340 $X2=1.2690 $Y2=0.2340
r19 77 79 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.5805 $Y=0.1350 $X2=1.5930 $Y2=0.1350
r20 76 77 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.5660 $Y=0.1350 $X2=1.5805 $Y2=0.1350
r21 74 76 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.5515 $Y=0.1350 $X2=1.5660 $Y2=0.1350
r22 73 74 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.5390 $Y=0.1350 $X2=1.5515 $Y2=0.1350
r23 71 73 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.5265 $Y=0.1350 $X2=1.5390 $Y2=0.1350
r24 70 71 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.5120 $Y=0.1350 $X2=1.5265 $Y2=0.1350
r25 68 70 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.4975 $Y=0.1350 $X2=1.5120 $Y2=0.1350
r26 67 68 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.4850 $Y=0.1350 $X2=1.4975 $Y2=0.1350
r27 65 67 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.4725 $Y=0.1350 $X2=1.4850 $Y2=0.1350
r28 64 65 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.4580 $Y=0.1350 $X2=1.4725 $Y2=0.1350
r29 62 64 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=1.4435 $Y=0.1350 $X2=1.4580 $Y2=0.1350
r30 60 62 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=1.4405 $Y=0.1350 $X2=1.4435 $Y2=0.1350
r31 59 60 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=1.4310
+ $Y=0.1350 $X2=1.4405 $Y2=0.1350
r32 2 59 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=1.4215
+ $Y=0.1350 $X2=1.4310 $Y2=0.1350
r33 29 55 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3770 $Y=0.2340 $X2=1.3770 $Y2=0.2125
r34 56 59 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.4310 $Y=0.1350
+ $X2=1.4310 $Y2=0.1350
r35 24 56 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.4040
+ $Y=0.1350 $X2=1.4310 $Y2=0.1350
r36 24 28 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.4040 $Y=0.1350 $X2=1.3770 $Y2=0.1350
r37 23 28 7.44771 $w=1.42162e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3770 $Y=0.1720 $X2=1.3770 $Y2=0.1350
r38 23 55 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=1.3770
+ $Y=0.1720 $X2=1.3770 $Y2=0.2125
r39 28 54 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.3770
+ $Y=0.1350 $X2=1.3770 $Y2=0.1125
r40 53 54 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.3770
+ $Y=0.0900 $X2=1.3770 $Y2=0.1125
r41 22 27 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3770 $Y=0.0630 $X2=1.3770 $Y2=0.0360
r42 22 53 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.3770
+ $Y=0.0630 $X2=1.3770 $Y2=0.0900
r43 52 51 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.1510 $Y=0.0675 $X2=1.1485 $Y2=0.0675
r44 50 51 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.1440 $Y=0.0675 $X2=1.1485 $Y2=0.0675
r45 6 50 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.1320 $Y=0.0675 $X2=1.1440 $Y2=0.0675
r46 16 6 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.1195 $Y=0.0675 $X2=1.1320 $Y2=0.0675
r47 49 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.1170 $Y=0.0675 $X2=1.1195 $Y2=0.0675
r48 27 47 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3770 $Y=0.0360 $X2=1.3500 $Y2=0.0360
r49 6 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.1340 $Y=0.0675
+ $X2=1.1340 $Y2=0.0360
r50 46 47 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=1.3095
+ $Y=0.0360 $X2=1.3500 $Y2=0.0360
r51 45 46 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=1.2850
+ $Y=0.0360 $X2=1.3095 $Y2=0.0360
r52 21 25 3.60008 $w=1.51951e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.2715 $Y=0.0360 $X2=1.2510 $Y2=0.0360
r53 21 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.2715
+ $Y=0.0360 $X2=1.2850 $Y2=0.0360
r54 42 43 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.1340
+ $Y=0.0360 $X2=1.1475 $Y2=0.0360
r55 40 43 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.0360 $X2=1.1475 $Y2=0.0360
r56 39 40 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.1880
+ $Y=0.0360 $X2=1.1610 $Y2=0.0360
r57 38 39 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.2150
+ $Y=0.0360 $X2=1.1880 $Y2=0.0360
r58 19 25 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.2330
+ $Y=0.0360 $X2=1.2510 $Y2=0.0360
r59 19 38 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.2330
+ $Y=0.0360 $X2=1.2150 $Y2=0.0360
r60 25 37 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.2510
+ $Y=0.0360 $X2=1.2510 $Y2=0.0540
r61 36 37 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.2510
+ $Y=0.0665 $X2=1.2510 $Y2=0.0540
r62 35 36 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.2510
+ $Y=0.0755 $X2=1.2510 $Y2=0.0665
r63 34 35 3.38125 $w=1.3e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=1.2510
+ $Y=0.0900 $X2=1.2510 $Y2=0.0755
r64 33 34 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.2510
+ $Y=0.1025 $X2=1.2510 $Y2=0.0900
r65 20 26 3.2503 $w=1.53684e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.2510 $Y=0.1160 $X2=1.2510 $Y2=0.1350
r66 20 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.2510
+ $Y=0.1160 $X2=1.2510 $Y2=0.1025
r67 26 31 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.2510
+ $Y=0.1350 $X2=1.2690 $Y2=0.1350
r68 11 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=1.2690
+ $Y=0.1350 $X2=1.2690 $Y2=0.1350
r69 1 31 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.2690 $Y=0.1350
+ $X2=1.2690 $Y2=0.1350
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%noxref_34 VSS 1
c1 1 VSS 0.0108217f
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%MH VSS 10 39 42 50 52 12 13 3 15 4 14 18 11 20 19
+ 17 1
c1 1 VSS 0.00342157f
c2 3 VSS 0.00674707f
c3 4 VSS 0.00346762f
c4 10 VSS 0.0793746f
c5 11 VSS 0.00225377f
c6 12 VSS 0.00216727f
c7 13 VSS 0.00233139f
c8 14 VSS 0.000465968f
c9 15 VSS 0.00031816f
c10 16 VSS 0.000201931f
c11 17 VSS 0.0111118f
c12 18 VSS 0.00278074f
c13 19 VSS 0.0002223f
c14 20 VSS 0.000130874f
c15 21 VSS 0.00196534f
c16 22 VSS 0.00287244f
r1 52 51 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.0675 $X2=0.7705 $Y2=0.0675
r2 12 51 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7580 $Y=0.0675 $X2=0.7705 $Y2=0.0675
r3 11 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.0675 $X2=0.7000 $Y2=0.0675
r4 50 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.0675 $X2=0.6875 $Y2=0.0675
r5 3 46 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7290 $Y=0.0675
+ $X2=0.7470 $Y2=0.0900
r6 46 47 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.7470
+ $Y=0.0900 $X2=0.7470 $Y2=0.1025
r7 45 47 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.7470
+ $Y=0.1135 $X2=0.7470 $Y2=0.1025
r8 44 45 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.7470
+ $Y=0.1425 $X2=0.7470 $Y2=0.1135
r9 43 44 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.7470
+ $Y=0.1655 $X2=0.7470 $Y2=0.1425
r10 14 19 3.01468 $w=1.741e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.7470
+ $Y=0.1780 $X2=0.7470 $Y2=0.1980
r11 14 43 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.7470
+ $Y=0.1780 $X2=0.7470 $Y2=0.1655
r12 19 37 1.73214 $w=1.61034e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7470 $Y=0.1980 $X2=0.7615 $Y2=0.1980
r13 42 41 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8270 $Y=0.2025 $X2=0.8245 $Y2=0.2025
r14 40 41 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8200 $Y=0.2025 $X2=0.8245 $Y2=0.2025
r15 4 40 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8080 $Y=0.2025 $X2=0.8200 $Y2=0.2025
r16 13 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.2025 $X2=0.8080 $Y2=0.2025
r17 39 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.2025 $X2=0.7955 $Y2=0.2025
r18 36 37 1.63233 $w=1.3e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.7685
+ $Y=0.1980 $X2=0.7615 $Y2=0.1980
r19 35 36 0.816164 $w=1.3e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.7720
+ $Y=0.1980 $X2=0.7685 $Y2=0.1980
r20 34 35 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1980 $X2=0.7720 $Y2=0.1980
r21 15 20 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7965 $Y=0.1980 $X2=0.8100 $Y2=0.1980
r22 15 34 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7965
+ $Y=0.1980 $X2=0.7830 $Y2=0.1980
r23 4 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8100 $Y=0.2025
+ $X2=0.8100 $Y2=0.2160
r24 16 21 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.2160 $X2=0.8100 $Y2=0.2340
r25 16 20 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.2160 $X2=0.8100 $Y2=0.1980
r26 21 33 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8100 $Y=0.2340 $X2=0.8235 $Y2=0.2340
r27 32 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.2340 $X2=0.8235 $Y2=0.2340
r28 31 32 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.2340 $X2=0.8370 $Y2=0.2340
r29 30 31 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.2340 $X2=0.8640 $Y2=0.2340
r30 17 22 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9180 $Y=0.2340 $X2=0.9450 $Y2=0.2340
r31 17 30 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.2340 $X2=0.8910 $Y2=0.2340
r32 22 29 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.2340 $X2=0.9450 $Y2=0.2125
r33 28 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1945 $X2=0.9450 $Y2=0.2125
r34 27 28 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1780 $X2=0.9450 $Y2=0.1945
r35 26 27 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1655 $X2=0.9450 $Y2=0.1780
r36 25 26 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1540 $X2=0.9450 $Y2=0.1655
r37 24 25 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1350 $X2=0.9450 $Y2=0.1540
r38 18 24 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1160 $X2=0.9450 $Y2=0.1350
r39 10 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.9450
+ $Y=0.1350 $X2=0.9450 $Y2=0.1350
r40 1 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.9450 $Y=0.1350
+ $X2=0.9450 $Y2=0.1350
r41 3 12 1e-05
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%PU1 VSS 12 13 24 8 2 7 1 9
c1 1 VSS 0.00471965f
c2 2 VSS 0.00468046f
c3 7 VSS 0.00218369f
c4 8 VSS 0.0021737f
c5 9 VSS 0.016649f
r1 24 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.2025 $X2=0.7705 $Y2=0.2025
r2 8 23 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7580 $Y=0.2025 $X2=0.7705 $Y2=0.2025
r3 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7560 $Y=0.2025
+ $X2=0.7560 $Y2=0.2340
r4 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7425
+ $Y=0.2340 $X2=0.7560 $Y2=0.2340
r5 19 20 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7245
+ $Y=0.2340 $X2=0.7425 $Y2=0.2340
r6 18 19 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7065
+ $Y=0.2340 $X2=0.7245 $Y2=0.2340
r7 17 18 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.2340 $X2=0.7065 $Y2=0.2340
r8 16 17 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6730
+ $Y=0.2340 $X2=0.6930 $Y2=0.2340
r9 15 16 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.6325
+ $Y=0.2340 $X2=0.6730 $Y2=0.2340
r10 14 15 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.2340 $X2=0.6325 $Y2=0.2340
r11 9 14 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5825
+ $Y=0.2340 $X2=0.5940 $Y2=0.2340
r12 1 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2025
+ $X2=0.5940 $Y2=0.2340
r13 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.2025 $X2=0.6085 $Y2=0.2025
r14 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.2025 $X2=0.6085 $Y2=0.2025
r15 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2025 $X2=0.5940 $Y2=0.2025
r16 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.2025 $X2=0.5795 $Y2=0.2025
r17 2 8 1e-05
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%SI VSS 14 3 9 12 8 4 1 6 5 10
c1 1 VSS 0.00312002f
c2 3 VSS 0.00687061f
c3 4 VSS 0.00153847f
c4 5 VSS 0.00159404f
c5 6 VSS 0.00171495f
c6 7 VSS 0.00173275f
c7 8 VSS 0.00717346f
c8 9 VSS 0.00167402f
c9 10 VSS 0.00162547f
c10 11 VSS 0.00353545f
c11 12 VSS 0.00158673f
r1 8 11 3.59766 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.7245
+ $Y=0.0360 $X2=0.7020 $Y2=0.0360
r2 7 12 2.45586 $w=1.44e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.0540 $X2=0.7020 $Y2=0.0665
r3 7 11 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.0540 $X2=0.7020 $Y2=0.0360
r4 12 19 1.40651 $w=1.51875e-08 $l=1.45774e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7020 $Y=0.0665 $X2=0.6885 $Y2=0.0720
r5 18 19 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.6730
+ $Y=0.0720 $X2=0.6885 $Y2=0.0720
r6 6 10 1.03257 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6595 $Y=0.0720 $X2=0.6480 $Y2=0.0720
r7 6 18 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6595
+ $Y=0.0720 $X2=0.6730 $Y2=0.0720
r8 5 17 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6480 $Y=0.0935 $X2=0.6480 $Y2=0.1150
r9 5 10 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6480 $Y=0.0935 $X2=0.6480 $Y2=0.0720
r10 16 17 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6345 $Y=0.1150 $X2=0.6480 $Y2=0.1150
r11 9 16 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.1150 $X2=0.6345 $Y2=0.1150
r12 14 4 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1250
r13 4 9 1.15159 $w=1.75e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1250 $X2=0.6210 $Y2=0.1150
r14 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1350
r15 14 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6210 $Y=0.1350
+ $X2=0.6210 $Y2=0.1350
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%NET54 VSS 15 34 35 37 11 2 13 10 1 12 3
c1 1 VSS 0.00606885f
c2 2 VSS 0.00605526f
c3 3 VSS 0.00344091f
c4 10 VSS 0.00448246f
c5 11 VSS 0.00333609f
c6 12 VSS 0.00266303f
c7 13 VSS 0.00530756f
r1 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.2025 $X2=0.6460 $Y2=0.2025
r2 37 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.2025 $X2=0.6335 $Y2=0.2025
r3 35 33 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r4 2 33 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5400 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r5 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.2025 $X2=0.5400 $Y2=0.2025
r6 34 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.2025 $X2=0.5255 $Y2=0.2025
r7 3 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.2025
+ $X2=0.6480 $Y2=0.1980
r8 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.2025
+ $X2=0.5400 $Y2=0.1980
r9 29 30 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6345
+ $Y=0.1980 $X2=0.6480 $Y2=0.1980
r10 28 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1980 $X2=0.6345 $Y2=0.1980
r11 27 28 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.6055
+ $Y=0.1980 $X2=0.6210 $Y2=0.1980
r12 26 27 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.5895
+ $Y=0.1980 $X2=0.6055 $Y2=0.1980
r13 25 26 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5780
+ $Y=0.1980 $X2=0.5895 $Y2=0.1980
r14 24 25 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1980 $X2=0.5780 $Y2=0.1980
r15 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5535
+ $Y=0.1980 $X2=0.5670 $Y2=0.1980
r16 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1980 $X2=0.5535 $Y2=0.1980
r17 21 22 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5265
+ $Y=0.1980 $X2=0.5400 $Y2=0.1980
r18 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1980 $X2=0.5265 $Y2=0.1980
r19 19 20 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.1980 $X2=0.5130 $Y2=0.1980
r20 18 19 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4635
+ $Y=0.1980 $X2=0.4860 $Y2=0.1980
r21 17 18 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4545
+ $Y=0.1980 $X2=0.4635 $Y2=0.1980
r22 16 17 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4455
+ $Y=0.1980 $X2=0.4545 $Y2=0.1980
r23 13 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.1980 $X2=0.4455 $Y2=0.1980
r24 1 13 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.1980
r25 15 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r26 10 14 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4340 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r27 1 10 1e-05
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%SE VSS 24 5 6 15 8 12 14 10 9 7 11 1 2 13
c1 1 VSS 0.0102872f
c2 2 VSS 0.0044705f
c3 5 VSS 0.0822689f
c4 6 VSS 0.0449104f
c5 7 VSS 0.00508101f
c6 8 VSS 0.00374249f
c7 9 VSS 0.00172117f
c8 10 VSS 0.0035058f
c9 11 VSS 0.00691719f
c10 12 VSS 0.00149892f
c11 13 VSS 0.00704062f
c12 14 VSS 0.00215183f
c13 15 VSS 0.00700341f
r1 2 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1350
+ $X2=0.5670 $Y2=0.1350
r2 6 2 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1350
r3 14 30 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.5670 $Y=0.0720 $X2=0.5670
+ $Y2=0.0810
r4 35 36 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1250 $X2=0.5670 $Y2=0.1350
r5 34 35 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1150 $X2=0.5670 $Y2=0.1250
r6 33 34 3.96423 $w=1.3e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0980 $X2=0.5670 $Y2=0.1150
r7 10 33 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0855 $X2=0.5670 $Y2=0.0980
r8 10 30 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.5670 $Y=0.0855 $X2=0.5670
+ $Y2=0.0810
r9 10 14 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.0855 $X2=0.5670 $Y2=0.0720
r10 29 30 37.7767 $w=1.3e-08 $l=1.62e-07 $layer=M2 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0810 $X2=0.5670 $Y2=0.0810
r11 28 29 37.7767 $w=1.3e-08 $l=1.62e-07 $layer=M2 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0810 $X2=0.4050 $Y2=0.0810
r12 15 28 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.2315
+ $Y=0.0810 $X2=0.2430 $Y2=0.0810
r13 8 12 10.3626 $w=1.39091e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.1845 $X2=0.2430 $Y2=0.1350
r14 8 13 10.3626 $w=1.39091e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.1845 $X2=0.2430 $Y2=0.2340
r15 25 26 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0810 $X2=0.2430 $Y2=0.1080
r16 25 28 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.2430 $Y=0.0810
+ $X2=0.2430 $Y2=0.0810
r17 7 25 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0585 $X2=0.2430 $Y2=0.0810
r18 7 11 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0585 $X2=0.2430 $Y2=0.0360
r19 12 26 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2430 $Y2=0.1080
r20 24 9 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2800
+ $Y=0.1350 $X2=0.2615 $Y2=0.1350
r21 9 12 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2615 $Y=0.1350 $X2=0.2430 $Y2=0.1350
r22 24 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2800 $Y=0.1350
+ $X2=0.2765 $Y2=0.1350
r23 20 22 4.72579 $w=1.53e-08 $l=8e-09 $layer=LIG $thickness=4.8e-08 $X=0.2845
+ $Y=0.1350 $X2=0.2765 $Y2=0.1350
r24 1 19 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.2880
+ $Y=0.1350 $X2=0.2980 $Y2=0.1350
r25 1 20 1.73797 $w=1.72143e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.2880 $Y=0.1350 $X2=0.2845 $Y2=0.1350
r26 5 19 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2980 $Y2=0.1350
r27 5 20 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2845 $Y2=0.1350
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%CLKN VSS 13 14 15 70 72 7 26 22 1 17 21 18 19 8
+ 28 20 16 23 2 24 3 25 27
c1 1 VSS 0.00379203f
c2 2 VSS 0.000155055f
c3 3 VSS 0.000111358f
c4 7 VSS 0.00871234f
c5 8 VSS 0.00878052f
c6 13 VSS 0.0801479f
c7 14 VSS 0.00436511f
c8 15 VSS 0.00444025f
c9 16 VSS 0.00818386f
c10 17 VSS 0.00820122f
c11 18 VSS 0.00406823f
c12 19 VSS 0.00610961f
c13 20 VSS 0.00692f
c14 21 VSS 0.00507157f
c15 22 VSS 0.00258491f
c16 23 VSS 0.000820943f
c17 24 VSS 0.00163847f
c18 25 VSS 0.00377858f
c19 26 VSS 0.00182756f
c20 27 VSS 0.00414354f
c21 28 VSS 0.0348042f
r1 72 71 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r2 17 71 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r3 70 69 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r4 16 69 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r5 8 67 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0550 $Y2=0.2340
r6 7 62 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0550 $Y2=0.0360
r7 66 67 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.2340 $X2=0.0550 $Y2=0.2340
r8 21 66 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0460 $Y2=0.2340
r9 21 27 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0180 $Y2=0.2340
r10 61 62 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.0360 $X2=0.0550 $Y2=0.0360
r11 20 61 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0460 $Y2=0.0360
r12 20 25 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0180 $Y2=0.0360
r13 27 58 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.2340 $X2=0.0180 $Y2=0.2125
r14 25 57 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0360 $X2=0.0180 $Y2=0.0540
r15 1 54 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1260
r16 13 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r17 19 26 9.39335 $w=1.38427e-08 $l=4.60245e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1630 $X2=0.0165 $Y2=0.1170
r18 19 58 11.5429 $w=1.3e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1630 $X2=0.0180 $Y2=0.2125
r19 56 57 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0720 $X2=0.0180 $Y2=0.0540
r20 18 26 3.9134 $w=1.47857e-08 $l=2.25499e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.0945 $X2=0.0165 $Y2=0.1170
r21 18 56 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0945 $X2=0.0180 $Y2=0.0720
r22 2 49 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7830 $Y=0.1350
+ $X2=0.7830 $Y2=0.1260
r23 14 2 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.7830
+ $Y=0.1350 $X2=0.7830 $Y2=0.1350
r24 22 54 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1055 $X2=0.1350 $Y2=0.1260
r25 51 52 1.90199 $w=1.38333e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.0255 $Y=0.1170 $X2=0.0345 $Y2=0.1170
r26 26 51 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0165
+ $Y=0.1170 $X2=0.0255 $Y2=0.1170
r27 23 49 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.0890 $X2=0.7830 $Y2=0.1260
r28 47 48 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1170 $X2=0.1595 $Y2=0.1170
r29 47 54 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1350 $Y=0.1170
+ $X2=0.1350 $Y2=0.1260
r30 46 47 11.8927 $w=1.3e-08 $l=5.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.0840
+ $Y=0.1170 $X2=0.1350 $Y2=0.1170
r31 45 46 11.8927 $w=1.3e-08 $l=5.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.0330
+ $Y=0.1170 $X2=0.0840 $Y2=0.1170
r32 45 52 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.0330 $Y=0.1170
+ $X2=0.0345 $Y2=0.1170
r33 43 48 9.91056 $w=1.3e-08 $l=4.25e-08 $layer=M2 $thickness=3.6e-08 $X=0.2020
+ $Y=0.1170 $X2=0.1595 $Y2=0.1170
r34 42 43 47.3375 $w=1.3e-08 $l=2.03e-07 $layer=M2 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1170 $X2=0.2020 $Y2=0.1170
r35 39 40 37.7767 $w=1.3e-08 $l=1.62e-07 $layer=M2 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1170 $X2=1.1070 $Y2=0.1170
r36 38 39 37.7767 $w=1.3e-08 $l=1.62e-07 $layer=M2 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1170 $X2=0.9450 $Y2=0.1170
r37 38 49 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.7830 $Y=0.1170
+ $X2=0.7830 $Y2=0.1260
r38 28 38 24.6015 $w=1.3e-08 $l=1.055e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.6775 $Y=0.1170 $X2=0.7830 $Y2=0.1170
r39 28 42 63.5442 $w=1.3e-08 $l=2.725e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.6775 $Y=0.1170 $X2=0.4050 $Y2=0.1170
r40 34 40 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=1.1070 $Y=0.1260
+ $X2=1.1070 $Y2=0.1170
r41 24 34 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.1070 $X2=1.1070 $Y2=0.1260
r42 15 3 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=1.1070
+ $Y=0.1350 $X2=1.1070 $Y2=0.1350
r43 3 34 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.1070 $Y=0.1350
+ $X2=1.1070 $Y2=0.1260
r44 8 17 1e-05
r45 7 16 1e-05
.ends

.subckt PM_SDFLx4_ASAP7_75t_R%CLKB VSS 15 16 17 18 78 80 10 9 29 27 22 21 1 28
+ 26 23 4 25 20 19 24 2 3
c1 1 VSS 9.38066e-20
c2 2 VSS 0.00010909f
c3 3 VSS 0.000109999f
c4 4 VSS 0.000253844f
c5 9 VSS 0.00785857f
c6 10 VSS 0.00847284f
c7 15 VSS 0.0051754f
c8 16 VSS 0.00433613f
c9 17 VSS 0.00466377f
c10 18 VSS 0.00533409f
c11 19 VSS 0.0104611f
c12 20 VSS 0.0105333f
c13 21 VSS 0.00706895f
c14 22 VSS 0.00374122f
c15 23 VSS 0.000350418f
c16 24 VSS 0.00168228f
c17 25 VSS 0.00134973f
c18 26 VSS 0.001842f
c19 27 VSS 0.00626526f
c20 28 VSS 0.00253519f
c21 29 VSS 0.0440796f
r1 19 9 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0675 $X2=0.1600 $Y2=0.0675
r2 80 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1475 $Y2=0.0675
r3 20 10 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1600 $Y2=0.2025
r4 78 20 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r5 9 73 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0675
+ $X2=0.1620 $Y2=0.0360
r6 15 69 2.79569 $w=1.27128e-07 $l=5e-10 $layer=LIG $thickness=5.21026e-08
+ $X=0.6750 $Y=0.1350 $X2=0.6745 $Y2=0.1350
r7 10 66 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r8 73 74 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r9 21 73 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1505
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r10 3 62 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.0530 $Y=0.1350
+ $X2=1.0530 $Y2=0.1440
r11 17 3 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=1.0530
+ $Y=0.1350 $X2=1.0530 $Y2=0.1350
r12 2 59 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8370 $Y=0.1350
+ $X2=0.8370 $Y2=0.1440
r13 16 2 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.8370
+ $Y=0.1350 $X2=0.8370 $Y2=0.1350
r14 69 70 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.6745
+ $Y=0.1350 $X2=0.6845 $Y2=0.1350
r15 1 70 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.6875 $Y=0.1350 $X2=0.6845 $Y2=0.1350
r16 1 72 5.02115 $w=1.53e-08 $l=8.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.6875
+ $Y=0.1350 $X2=0.6960 $Y2=0.1350
r17 66 67 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r18 27 54 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2340 $X2=0.1890 $Y2=0.2125
r19 27 67 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2340 $X2=0.1755 $Y2=0.2340
r20 28 53 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.1890 $Y2=0.0540
r21 28 74 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1755 $Y2=0.0360
r22 25 62 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1160 $X2=1.0530 $Y2=0.1440
r23 24 59 10.7267 $w=1.3e-08 $l=4.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.0980 $X2=0.8370 $Y2=0.1440
r24 55 72 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6930 $Y=0.1440
+ $X2=0.6960 $Y2=0.1350
r25 23 55 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1250 $X2=0.6930 $Y2=0.1440
r26 52 53 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0720 $X2=0.1890 $Y2=0.0540
r27 51 52 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0920 $X2=0.1890 $Y2=0.0720
r28 50 54 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1810 $X2=0.1890 $Y2=0.2125
r29 49 50 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1530 $X2=0.1890 $Y2=0.1810
r30 22 49 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1235 $X2=0.1890 $Y2=0.1530
r31 22 51 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1235 $X2=0.1890 $Y2=0.0920
r32 47 48 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M2 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1530 $X2=1.0915 $Y2=0.1530
r33 47 62 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=1.0530 $Y=0.1530
+ $X2=1.0530 $Y2=0.1440
r34 46 47 25.1845 $w=1.3e-08 $l=1.08e-07 $layer=M2 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1530 $X2=1.0530 $Y2=0.1530
r35 45 46 25.1845 $w=1.3e-08 $l=1.08e-07 $layer=M2 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1530 $X2=0.9450 $Y2=0.1530
r36 45 59 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.8370 $Y=0.1530
+ $X2=0.8370 $Y2=0.1440
r37 44 45 16.7897 $w=1.3e-08 $l=7.2e-08 $layer=M2 $thickness=3.6e-08 $X=0.7650
+ $Y=0.1530 $X2=0.8370 $Y2=0.1530
r38 43 44 16.7897 $w=1.3e-08 $l=7.2e-08 $layer=M2 $thickness=3.6e-08 $X=0.6930
+ $Y=0.1530 $X2=0.7650 $Y2=0.1530
r39 43 55 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.6930 $Y=0.1530
+ $X2=0.6930 $Y2=0.1440
r40 42 43 58.7638 $w=1.3e-08 $l=2.52e-07 $layer=M2 $thickness=3.6e-08 $X=0.4410
+ $Y=0.1530 $X2=0.6930 $Y2=0.1530
r41 41 42 58.7638 $w=1.3e-08 $l=2.52e-07 $layer=M2 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1530 $X2=0.4410 $Y2=0.1530
r42 41 49 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1890 $Y=0.1530
+ $X2=0.1890 $Y2=0.1530
r43 29 38 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=1.1365
+ $Y=0.1530 $X2=1.1610 $Y2=0.1530
r44 29 48 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M2 $thickness=3.6e-08 $X=1.1365
+ $Y=0.1530 $X2=1.0915 $Y2=0.1530
r45 35 38 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=1.1610 $Y=0.1440
+ $X2=1.1610 $Y2=0.1530
r46 26 35 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.1610
+ $Y=0.1160 $X2=1.1610 $Y2=0.1440
r47 18 4 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=1.1610
+ $Y=0.1350 $X2=1.1610 $Y2=0.1350
r48 4 35 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.1610 $Y=0.1350
+ $X2=1.1610 $Y2=0.1440
.ends


*
.SUBCKT SDFLx4_ASAP7_75t_R VSS VDD CLK SE D SI QN
*
* VSS VSS
* VDD VDD
* CLK CLK
* SE SE
* D D
* SI SI
* QN QN
*
*

MM20 N_MM20_d N_MM20_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM23 N_MM23_d N_MM23_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM30 N_MM30_d N_MM31_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM29 N_MM29_d N_MM26_g N_MM29_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM28 N_MM28_d N_MM0_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM27 N_MM27_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM2_g N_MM5_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM1_g N_MM9_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM6_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM12 N_MM12_d N_MM12_g N_MM12_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM17 N_MM17_d N_MM17_g N_MM17_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM16 N_MM16_d N_MM16_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM14 N_MM14_d N_MM14_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24 N_MM24_d N_MM24_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@4 N_MM24@4_d N_MM24@4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@3 N_MM24@3_d N_MM24@3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@2 N_MM24@2_d N_MM24@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM21 N_MM21_d N_MM20_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM22 N_MM22_d N_MM23_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM31 N_MM31_d N_MM31_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM26 N_MM26_d N_MM26_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g N_MM3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g N_MM2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM6_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM13 N_MM13_d N_MM13_g N_MM13_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM18 N_MM18_d N_MM12_g N_MM18_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM19 N_MM19_d N_MM16_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM15 N_MM15_d N_MM14_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25 N_MM25_d N_MM24_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@4 N_MM25@4_d N_MM24@4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@3 N_MM25@3_d N_MM24@3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@2 N_MM25@2_d N_MM24@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "SDFLx4_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "SDFLx4_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_SDFLx4_ASAP7_75t_R%NET066 VSS N_MM29_s N_MM28_d N_NET066_1
+ PM_SDFLx4_ASAP7_75t_R%NET066
cc_1 N_NET066_1 N_MM26_g 0.0172893f
cc_2 N_NET066_1 N_MM0_g 0.0172791f
x_PM_SDFLx4_ASAP7_75t_R%NET067 VSS N_MM27_d N_MM5_s N_NET067_1
+ PM_SDFLx4_ASAP7_75t_R%NET067
cc_3 N_NET067_1 N_MM3_g 0.0173965f
cc_4 N_NET067_1 N_MM2_g 0.0172782f
x_PM_SDFLx4_ASAP7_75t_R%noxref_31 VSS N_noxref_31_1
+ PM_SDFLx4_ASAP7_75t_R%noxref_31
cc_5 N_noxref_31_1 N_MM31_g 0.00134383f
cc_6 N_noxref_31_1 N_SEN_11 0.0376926f
cc_7 N_noxref_31_1 N_noxref_30_1 0.00122999f
x_PM_SDFLx4_ASAP7_75t_R%noxref_32 VSS N_noxref_32_1
+ PM_SDFLx4_ASAP7_75t_R%noxref_32
cc_8 N_noxref_32_1 N_MM26_g 0.0015056f
cc_9 N_noxref_32_1 N_SEN_10 0.000921353f
cc_10 N_noxref_32_1 N_PD1_7 0.0354762f
cc_11 N_noxref_32_1 N_noxref_30_1 0.00766401f
x_PM_SDFLx4_ASAP7_75t_R%noxref_30 VSS N_noxref_30_1
+ PM_SDFLx4_ASAP7_75t_R%noxref_30
cc_12 N_noxref_30_1 N_MM31_g 0.00134084f
cc_13 N_noxref_30_1 N_SEN_10 0.0378271f
x_PM_SDFLx4_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_SDFLx4_ASAP7_75t_R%noxref_24
cc_14 N_noxref_24_1 N_MM20_g 0.00144599f
cc_15 N_noxref_24_1 N_CLKN_25 5.64802e-20
cc_16 N_noxref_24_1 N_CLKN_26 6.89282e-20
cc_17 N_noxref_24_1 N_CLKN_8 7.44569e-20
cc_18 N_noxref_24_1 N_CLKN_17 9.04359e-20
cc_19 N_noxref_24_1 N_CLKN_19 0.000125558f
cc_20 N_noxref_24_1 N_CLKN_18 0.00017473f
cc_21 N_noxref_24_1 N_CLKN_7 0.000501466f
cc_22 N_noxref_24_1 N_CLKN_16 0.0374348f
x_PM_SDFLx4_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_SDFLx4_ASAP7_75t_R%noxref_25
cc_23 N_noxref_25_1 N_MM20_g 0.0014493f
cc_24 N_noxref_25_1 N_CLKN_18 5.45523e-20
cc_25 N_noxref_25_1 N_CLKN_27 5.78818e-20
cc_26 N_noxref_25_1 N_CLKN_7 7.33354e-20
cc_27 N_noxref_25_1 N_CLKN_16 8.98865e-20
cc_28 N_noxref_25_1 N_CLKN_19 0.000268357f
cc_29 N_noxref_25_1 N_CLKN_8 0.000502373f
cc_30 N_noxref_25_1 N_CLKN_17 0.0374213f
cc_31 N_noxref_25_1 N_noxref_24_1 0.00175947f
x_PM_SDFLx4_ASAP7_75t_R%PD5 VSS N_MM17_s N_MM16_d N_PD5_1
+ PM_SDFLx4_ASAP7_75t_R%PD5
cc_32 N_PD5_1 N_MM17_g 0.0170138f
cc_33 N_PD5_1 N_MM16_g 0.0170874f
x_PM_SDFLx4_ASAP7_75t_R%PD3 VSS N_MM9_s N_MM8_d N_PD3_4 N_PD3_5 N_PD3_1
+ PM_SDFLx4_ASAP7_75t_R%PD3
cc_34 N_PD3_4 N_CLKN_2 0.000828907f
cc_35 N_PD3_4 N_CLKN_23 0.000529847f
cc_36 N_PD3_4 N_MM1_g 0.0344404f
cc_37 N_PD3_4 N_CLKB_2 0.00197068f
cc_38 N_PD3_4 N_CLKB_24 0.00107607f
cc_39 N_PD3_4 N_MM10_g 0.0740804f
cc_40 N_PD3_5 N_MM11_g 0.0365879f
cc_41 N_PD3_1 N_MH_3 0.00120038f
cc_42 N_PD3_1 N_MH_12 0.00286077f
x_PM_SDFLx4_ASAP7_75t_R%noxref_27 VSS N_noxref_27_1
+ PM_SDFLx4_ASAP7_75t_R%noxref_27
cc_43 N_noxref_27_1 N_MM23_g 0.00135799f
cc_44 N_noxref_27_1 N_CLKB_19 7.44805e-20
cc_45 N_noxref_27_1 N_CLKB_22 0.0001133f
cc_46 N_noxref_27_1 N_CLKB_10 0.000416483f
cc_47 N_noxref_27_1 N_CLKB_20 0.037086f
cc_48 N_noxref_27_1 N_noxref_26_1 0.00123781f
x_PM_SDFLx4_ASAP7_75t_R%noxref_26 VSS N_noxref_26_1
+ PM_SDFLx4_ASAP7_75t_R%noxref_26
cc_49 N_noxref_26_1 N_MM23_g 0.00135654f
cc_50 N_noxref_26_1 N_CLKB_20 7.26656e-20
cc_51 N_noxref_26_1 N_CLKB_22 0.000112709f
cc_52 N_noxref_26_1 N_CLKB_9 0.00041704f
cc_53 N_noxref_26_1 N_CLKB_19 0.0371638f
x_PM_SDFLx4_ASAP7_75t_R%noxref_29 VSS N_noxref_29_1
+ PM_SDFLx4_ASAP7_75t_R%noxref_29
cc_54 N_noxref_29_1 N_MM31_g 0.00179604f
cc_55 N_noxref_29_1 N_CLKB_22 8.59806e-20
cc_56 N_noxref_29_1 N_CLKB_10 0.000136388f
cc_57 N_noxref_29_1 N_CLKB_20 0.000583831f
cc_58 N_noxref_29_1 N_noxref_27_1 0.00765313f
cc_59 N_noxref_29_1 N_noxref_28_1 0.00122493f
x_PM_SDFLx4_ASAP7_75t_R%PD2 VSS N_MM10_s N_MM11_d N_PD2_3 N_PD2_1
+ PM_SDFLx4_ASAP7_75t_R%PD2
cc_60 N_PD2_3 N_CLKB_2 0.000869035f
cc_61 N_PD2_3 N_CLKB_24 0.000209508f
cc_62 N_PD2_3 N_MM10_g 0.0334648f
cc_63 N_PD2_3 N_MM11_g 0.0345939f
cc_64 N_PD2_1 N_MH_13 0.000567901f
cc_65 N_PD2_1 N_MH_17 0.000672899f
cc_66 N_PD2_1 N_MH_4 0.00423497f
x_PM_SDFLx4_ASAP7_75t_R%noxref_28 VSS N_noxref_28_1
+ PM_SDFLx4_ASAP7_75t_R%noxref_28
cc_67 N_noxref_28_1 N_MM31_g 0.00179734f
cc_68 N_noxref_28_1 N_CLKB_22 8.55922e-20
cc_69 N_noxref_28_1 N_CLKB_9 0.000132949f
cc_70 N_noxref_28_1 N_CLKB_19 0.000586295f
cc_71 N_noxref_28_1 N_noxref_26_1 0.00765071f
x_PM_SDFLx4_ASAP7_75t_R%noxref_35 VSS N_noxref_35_1
+ PM_SDFLx4_ASAP7_75t_R%noxref_35
cc_72 N_noxref_35_1 N_MM13_g 0.0100532f
cc_73 N_noxref_35_1 N_MS_5 0.00089487f
cc_74 N_noxref_35_1 N_MS_3 0.00141174f
cc_75 N_noxref_35_1 N_MS_4 0.00211544f
cc_76 N_noxref_35_1 N_MS_12 0.0163877f
cc_77 N_noxref_35_1 N_MS_15 0.0163842f
cc_78 N_noxref_35_1 N_MS_14 0.0784683f
cc_79 N_noxref_35_1 N_MM6_g 0.00325555f
x_PM_SDFLx4_ASAP7_75t_R%CLK VSS CLK N_MM20_g N_CLK_4 N_CLK_5 N_CLK_1
+ PM_SDFLx4_ASAP7_75t_R%CLK
x_PM_SDFLx4_ASAP7_75t_R%PD1 VSS N_MM29_d N_MM5_d N_MM4_s N_PD1_9 N_PD1_7
+ N_PD1_1 N_PD1_8 N_PD1_2 PM_SDFLx4_ASAP7_75t_R%PD1
cc_80 N_PD1_9 N_SE_10 0.000494728f
cc_81 N_PD1_9 N_MM3_g 0.000236927f
cc_82 N_PD1_9 N_SE_15 0.000915413f
cc_83 N_PD1_9 N_SE_14 0.00602368f
cc_84 N_PD1_7 N_D_1 0.000791057f
cc_85 N_PD1_1 N_MM26_g 0.00172482f
cc_86 N_PD1_7 N_MM26_g 0.0352082f
cc_87 N_PD1_9 N_MM0_g 0.000241686f
cc_88 N_PD1_1 N_SEN_14 0.00183241f
cc_89 N_PD1_9 N_SEN_14 0.00454592f
cc_90 N_PD1_9 N_SEN_19 0.00669315f
cc_91 N_PD1_8 N_SI_5 0.000349179f
cc_92 N_PD1_2 N_SI_10 0.000382452f
cc_93 N_PD1_8 N_SI_1 0.000670662f
cc_94 N_PD1_9 N_SI_6 0.000750607f
cc_95 N_PD1_9 N_SI_10 0.00119487f
cc_96 N_PD1_9 N_SI_9 0.00190779f
cc_97 N_PD1_2 N_MM2_g 0.00195929f
cc_98 N_PD1_8 N_MM2_g 0.0351137f
cc_99 N_PD1_8 N_CLKB_29 0.000134964f
cc_100 N_PD1_8 N_CLKB_1 0.000745488f
cc_101 N_PD1_2 N_MM4_g 0.000776563f
cc_102 N_PD1_8 N_MM4_g 0.0334522f
cc_103 N_PD1_8 N_MH_11 0.000556474f
cc_104 N_PD1_2 N_MH_3 0.00116416f
cc_105 N_PD1_8 N_MH_3 0.00216804f
x_PM_SDFLx4_ASAP7_75t_R%noxref_33 VSS N_noxref_33_1
+ PM_SDFLx4_ASAP7_75t_R%noxref_33
cc_106 N_noxref_33_1 N_MM26_g 0.00162388f
cc_107 N_noxref_33_1 N_SEN_11 0.000815384f
cc_108 N_noxref_33_1 N_NET54_10 0.0355807f
cc_109 N_noxref_33_1 N_noxref_31_1 0.00764761f
cc_110 N_noxref_33_1 N_noxref_32_1 0.00123858f
x_PM_SDFLx4_ASAP7_75t_R%D VSS D N_MM26_g N_D_7 N_D_1 N_D_10 N_D_8 N_D_9 N_D_5
+ N_D_4 N_D_6 PM_SDFLx4_ASAP7_75t_R%D
cc_111 N_D_7 N_CLKN_28 0.00246055f
x_PM_SDFLx4_ASAP7_75t_R%SEN VSS N_MM0_g N_MM30_d N_MM31_d N_SEN_10 N_SEN_17
+ N_SEN_16 N_SEN_11 N_SEN_4 N_SEN_1 N_SEN_19 N_SEN_3 N_SEN_13 N_SEN_15 N_SEN_14
+ PM_SDFLx4_ASAP7_75t_R%SEN
cc_112 N_SEN_10 N_SE_11 0.000152069f
cc_113 N_SEN_10 N_SE_15 0.000741351f
cc_114 N_SEN_17 N_SE_8 0.000339253f
cc_115 N_SEN_16 N_SE_7 0.000340564f
cc_116 N_SEN_11 N_MM31_g 0.0157721f
cc_117 N_SEN_4 N_SE_1 0.000590857f
cc_118 N_SEN_1 N_SE_2 0.00158341f
cc_119 N_SEN_19 N_SE_14 0.000771116f
cc_120 N_SEN_17 N_SE_13 0.000797884f
cc_121 N_SEN_16 N_SE_11 0.00108138f
cc_122 N_SEN_4 N_MM31_g 0.00109982f
cc_123 N_SEN_3 N_MM31_g 0.00112029f
cc_124 N_SEN_13 N_SE_9 0.00198368f
cc_125 N_SEN_11 N_SE_1 0.00204775f
cc_126 N_SEN_15 N_SE_10 0.00305638f
cc_127 N_MM0_g N_MM3_g 0.00328047f
cc_128 N_SEN_14 N_SE_15 0.00420538f
cc_129 N_SEN_10 N_MM31_g 0.0544058f
cc_130 N_SEN_1 N_D_1 0.00218614f
cc_131 N_SEN_14 N_D_10 0.00121398f
cc_132 N_SEN_13 N_D_8 0.00132907f
cc_133 N_SEN_17 N_D_9 0.00170046f
cc_134 N_SEN_15 N_D_7 0.00192096f
cc_135 N_MM0_g N_MM26_g 0.00499653f
cc_136 N_SEN_14 N_D_5 0.00647049f
cc_137 N_SEN_13 N_D_4 0.00879584f
x_PM_SDFLx4_ASAP7_75t_R%noxref_36 VSS N_noxref_36_1
+ PM_SDFLx4_ASAP7_75t_R%noxref_36
cc_138 N_noxref_36_1 N_SS_3 0.00145621f
cc_139 N_noxref_36_1 N_SS_10 0.0374735f
cc_140 N_noxref_36_1 N_MM14_g 0.00152747f
x_PM_SDFLx4_ASAP7_75t_R%noxref_38 VSS N_noxref_38_1
+ PM_SDFLx4_ASAP7_75t_R%noxref_38
cc_141 N_noxref_38_1 N_SS_10 0.00110149f
cc_142 N_noxref_38_1 N_MM24_g 0.00176286f
cc_143 N_noxref_38_1 N_noxref_36_1 0.00753653f
x_PM_SDFLx4_ASAP7_75t_R%noxref_39 VSS N_noxref_39_1
+ PM_SDFLx4_ASAP7_75t_R%noxref_39
cc_144 N_noxref_39_1 N_SS_11 0.000808725f
cc_145 N_noxref_39_1 N_MM24_g 0.00180903f
cc_146 N_noxref_39_1 N_noxref_37_1 0.00766121f
cc_147 N_noxref_39_1 N_noxref_38_1 0.00124117f
x_PM_SDFLx4_ASAP7_75t_R%noxref_37 VSS N_noxref_37_1
+ PM_SDFLx4_ASAP7_75t_R%noxref_37
cc_148 N_noxref_37_1 N_SS_11 0.0377243f
cc_149 N_noxref_37_1 N_MM14_g 0.00167977f
cc_150 N_noxref_37_1 N_noxref_36_1 0.00121773f
x_PM_SDFLx4_ASAP7_75t_R%noxref_40 VSS N_noxref_40_1
+ PM_SDFLx4_ASAP7_75t_R%noxref_40
cc_151 N_noxref_40_1 N_MM24@2_g 0.00147423f
cc_152 N_noxref_40_1 N_QN_14 0.000832742f
x_PM_SDFLx4_ASAP7_75t_R%noxref_41 VSS N_noxref_41_1
+ PM_SDFLx4_ASAP7_75t_R%noxref_41
cc_153 N_noxref_41_1 N_MM24@2_g 0.00146661f
cc_154 N_noxref_41_1 N_QN_16 0.00083254f
cc_155 N_noxref_41_1 N_noxref_40_1 0.00177139f
x_PM_SDFLx4_ASAP7_75t_R%PD4 VSS N_MM18_s N_MM19_d N_PD4_4 N_PD4_5 N_PD4_1
+ PM_SDFLx4_ASAP7_75t_R%PD4
cc_156 N_PD4_4 N_CLKN_24 0.000205166f
cc_157 N_PD4_4 N_CLKN_3 0.000694533f
cc_158 N_PD4_4 N_MM12_g 0.0342012f
cc_159 N_PD4_4 N_CLKB_4 0.00225619f
cc_160 N_PD4_4 N_CLKB_26 0.000995754f
cc_161 N_PD4_4 N_MM17_g 0.0737343f
cc_162 N_PD4_5 N_SS_1 0.000812344f
cc_163 N_PD4_5 N_MM16_g 0.0351092f
cc_164 N_PD4_1 N_SH_5 0.00135725f
cc_165 N_PD4_1 N_SH_17 0.00115519f
cc_166 N_PD4_1 N_SH_18 0.00447389f
x_PM_SDFLx4_ASAP7_75t_R%QN VSS QN N_MM24_d N_MM24@4_d N_MM24@3_d N_MM24@2_d
+ N_MM25_d N_MM25@4_d N_MM25@3_d N_MM25@2_d N_QN_14 N_QN_16 N_QN_15 N_QN_13
+ N_QN_18 N_QN_17 N_QN_2 N_QN_3 N_QN_4 N_QN_1 PM_SDFLx4_ASAP7_75t_R%QN
cc_167 N_QN_14 N_SH_27 0.000154134f
cc_168 N_QN_14 N_SH_29 0.000162518f
cc_169 N_QN_14 N_MM24_g 0.00036064f
cc_170 N_QN_14 N_SH_22 0.000443759f
cc_171 N_QN_14 N_SH_23 0.000447028f
cc_172 N_QN_14 N_SH_2 0.00123431f
cc_173 N_QN_16 N_MM24@3_g 0.030554f
cc_174 N_QN_15 N_MM24_g 0.0305208f
cc_175 N_QN_13 N_MM24_g 0.0672424f
cc_176 N_QN_18 N_MM24@3_g 0.000905735f
cc_177 N_QN_17 N_MM24@3_g 0.000940826f
cc_178 N_QN_2 N_SH_24 0.0010025f
cc_179 N_QN_3 N_MM24@3_g 0.00176832f
cc_180 N_QN_4 N_MM24@3_g 0.00182086f
cc_181 N_QN_1 N_MM24_g 0.00208985f
cc_182 N_QN_2 N_MM24_g 0.00213306f
cc_183 N_QN_15 N_SH_2 0.00972167f
cc_184 N_QN_14 N_MM24@2_g 0.0367244f
cc_185 N_QN_13 N_MM24@4_g 0.0367778f
cc_186 N_QN_14 N_MM24@3_g 0.067686f
x_PM_SDFLx4_ASAP7_75t_R%SS VSS N_MM16_g N_MM15_d N_MM14_d N_SS_1 N_SS_12
+ N_SS_10 N_SS_11 N_SS_3 N_SS_14 N_SS_4 N_SS_17 N_SS_16 N_SS_13 N_SS_15
+ PM_SDFLx4_ASAP7_75t_R%SS
cc_187 N_MM16_g N_CLKB_26 0.000766302f
cc_188 N_MM16_g N_CLKB_29 0.000432307f
cc_189 N_SS_1 N_CLKB_4 0.00230703f
cc_190 N_SS_12 N_CLKB_26 0.00322949f
cc_191 N_MM16_g N_MM17_g 0.005109f
x_PM_SDFLx4_ASAP7_75t_R%MS VSS N_MM11_g N_MM6_d N_MM12_d N_MM7_d N_MM13_d
+ N_MS_13 N_MS_17 N_MS_4 N_MS_16 N_MS_15 N_MS_1 N_MS_5 N_MS_3 N_MS_12 N_MS_14
+ PM_SDFLx4_ASAP7_75t_R%MS
cc_192 N_MS_13 N_CLKN_3 0.000921599f
cc_193 N_MS_13 N_MM1_g 7.85539e-20
cc_194 N_MS_13 N_CLKN_28 0.000230468f
cc_195 N_MS_13 N_CLKN_24 0.00070555f
cc_196 N_MS_17 N_CLKN_28 0.000737717f
cc_197 N_MS_4 N_MM12_g 0.00159577f
cc_198 N_MS_16 N_CLKN_28 0.00245737f
cc_199 N_MS_13 N_MM12_g 0.0346047f
cc_200 N_MS_15 N_MM17_g 5.17217e-20
cc_201 N_MS_15 N_CLKB_25 0.000114133f
cc_202 N_MS_15 N_CLKB_24 0.000541504f
cc_203 N_MS_15 N_CLKB_29 0.000273273f
cc_204 N_MS_15 N_CLKB_2 0.000755831f
cc_205 N_MS_13 N_MM13_g 0.0175788f
cc_206 N_MS_16 N_CLKB_29 0.000882597f
cc_207 N_MS_1 N_CLKB_2 0.000902485f
cc_208 N_MS_4 N_CLKB_3 0.00370708f
cc_209 N_MS_5 N_MM13_g 0.00147576f
cc_210 N_MS_3 N_CLKB_3 0.00150024f
cc_211 N_MS_5 N_CLKB_25 0.00168157f
cc_212 N_MM11_g N_MM10_g 0.0033041f
cc_213 N_MS_16 N_CLKB_24 0.00361074f
cc_214 N_MS_4 N_MM13_g 0.00463078f
cc_215 N_MS_15 N_MM13_g 0.0552236f
x_PM_SDFLx4_ASAP7_75t_R%SH VSS N_MM14_g N_MM24_g N_MM24@4_g N_MM24@3_g
+ N_MM24@2_g N_MM12_s N_MM17_d N_MM13_s N_MM18_d N_SH_16 N_SH_6 N_SH_18 N_SH_17
+ N_SH_5 N_SH_19 N_SH_26 N_SH_20 N_SH_2 N_SH_24 N_SH_1 N_SH_28 N_SH_23 N_SH_21
+ N_SH_22 N_SH_27 N_SH_29 PM_SDFLx4_ASAP7_75t_R%SH
cc_216 N_SH_16 N_CLKN_24 8.80643e-20
cc_217 N_SH_6 N_CLKN_24 0.00199244f
cc_218 N_SH_18 N_CLKN_24 0.000330891f
cc_219 N_SH_18 N_CLKN_28 0.000386099f
cc_220 N_SH_17 N_MM12_g 0.0155755f
cc_221 N_SH_5 N_CLKN_3 0.000423625f
cc_222 N_SH_5 N_MM12_g 0.000981121f
cc_223 N_SH_19 N_CLKN_24 0.00102719f
cc_224 N_SH_6 N_MM12_g 0.00128879f
cc_225 N_SH_17 N_CLKN_3 0.00135155f
cc_226 N_SH_16 N_MM12_g 0.0537727f
cc_227 N_SH_16 N_CLKB_26 5.24639e-20
cc_228 N_SH_16 N_CLKB_25 6.52414e-20
cc_229 N_SH_18 N_CLKB_26 0.0028278f
cc_230 N_SH_26 N_CLKB_26 0.000160244f
cc_231 N_SH_5 N_CLKB_25 0.00155812f
cc_232 N_SH_20 N_CLKB_26 0.000207034f
cc_233 N_SH_5 N_CLKB_3 0.000222946f
cc_234 N_SH_6 N_CLKB_4 0.000332798f
cc_235 N_SH_17 N_MM13_g 0.0345578f
cc_236 N_SH_19 N_CLKB_26 0.000615331f
cc_237 N_SH_17 N_CLKB_3 0.000706157f
cc_238 N_SH_16 N_CLKB_4 0.000862353f
cc_239 N_SH_18 N_CLKB_29 0.000960642f
cc_240 N_SH_5 N_MM13_g 0.00132631f
cc_241 N_SH_6 N_MM17_g 0.00137626f
cc_242 N_SH_6 N_CLKB_26 0.00193944f
cc_243 N_SH_16 N_MM17_g 0.035436f
cc_244 N_SH_18 N_MS_4 0.000172521f
cc_245 N_SH_5 N_MS_4 0.000180201f
cc_246 N_SH_19 N_MS_4 0.000193581f
cc_247 N_SH_6 N_MS_4 0.00142271f
cc_248 N_SH_17 N_MS_4 0.000571315f
cc_249 N_SH_17 N_MS_15 0.000614991f
cc_250 N_SH_16 N_MS_13 0.000616334f
cc_251 N_SH_5 N_MS_5 0.00126096f
cc_252 N_SH_17 N_MS_5 0.00150569f
cc_253 N_SH_16 N_MS_4 0.00241456f
cc_254 N_SH_16 N_SS_10 9.15269e-20
cc_255 N_SH_2 N_SS_10 9.54403e-20
cc_256 N_SH_24 N_SS_10 0.000152189f
cc_257 N_SH_6 N_SS_10 0.000228342f
cc_258 N_SH_18 N_SS_10 0.000440877f
cc_259 N_SH_19 N_SS_10 0.000442266f
cc_260 N_MM14_g N_SS_11 0.0158137f
cc_261 N_SH_1 N_SS_1 0.000591203f
cc_262 N_SH_26 N_SS_1 0.000631315f
cc_263 N_SH_20 N_SS_3 0.000695555f
cc_264 N_SH_28 N_SS_14 0.000743323f
cc_265 N_SH_1 N_SS_4 0.0012544f
cc_266 N_SH_18 N_SS_17 0.00140842f
cc_267 N_SH_23 N_SS_17 0.00150946f
cc_268 N_MM14_g N_SS_4 0.00170784f
cc_269 N_MM14_g N_MM16_g 0.00192283f
cc_270 N_SH_21 N_SS_16 0.00201129f
cc_271 N_SH_1 N_SS_11 0.00215211f
cc_272 N_MM14_g N_SS_3 0.00244116f
cc_273 N_SH_22 N_SS_16 0.00248973f
cc_274 N_SH_20 N_SS_12 0.00272762f
cc_275 N_SH_26 N_SS_14 0.00319257f
cc_276 N_SH_26 N_SS_16 0.00325462f
cc_277 N_SH_18 N_SS_13 0.00329491f
cc_278 N_SH_26 N_SS_12 0.00426692f
cc_279 N_SH_18 N_SS_15 0.00556963f
cc_280 N_MM14_g N_SS_10 0.0557687f
x_PM_SDFLx4_ASAP7_75t_R%noxref_34 VSS N_noxref_34_1
+ PM_SDFLx4_ASAP7_75t_R%noxref_34
cc_281 N_noxref_34_1 N_MM1_g 0.00347922f
cc_282 N_noxref_34_1 N_MM4_g 0.00507027f
cc_283 N_noxref_34_1 N_CLKB_1 0.0068344f
cc_284 N_noxref_34_1 N_MH_3 0.00112726f
cc_285 N_noxref_34_1 N_MH_12 0.0166117f
cc_286 N_noxref_34_1 N_MH_11 0.0564589f
cc_287 N_noxref_34_1 N_PU1_8 0.0368025f
x_PM_SDFLx4_ASAP7_75t_R%MH VSS N_MM6_g N_MM1_d N_MM10_d N_MM4_d N_MM9_d N_MH_12
+ N_MH_13 N_MH_3 N_MH_15 N_MH_4 N_MH_14 N_MH_18 N_MH_11 N_MH_20 N_MH_19 N_MH_17
+ N_MH_1 PM_SDFLx4_ASAP7_75t_R%MH
cc_288 N_MH_12 N_CLKN_23 0.00102557f
cc_289 N_MH_13 N_MM1_g 0.015561f
cc_290 N_MH_3 N_CLKN_28 0.000482007f
cc_291 N_MH_15 N_CLKN_23 0.000771165f
cc_292 N_MH_4 N_MM1_g 0.0009002f
cc_293 N_MH_14 N_CLKN_2 0.000962488f
cc_294 N_MH_3 N_MM1_g 0.00117926f
cc_295 N_MH_13 N_CLKN_2 0.0016127f
cc_296 N_MH_18 N_CLKN_28 0.00165168f
cc_297 N_MH_14 N_CLKN_23 0.00827318f
cc_298 N_MH_12 N_MM1_g 0.05345f
cc_299 N_MH_3 N_SI_6 0.000372599f
cc_300 N_MH_14 N_SI_8 0.00149815f
cc_301 N_MH_3 N_SI_12 0.00179107f
cc_302 N_MH_14 N_SI_12 0.00327816f
cc_303 N_MH_11 N_MM13_g 4.39956e-20
cc_304 N_MH_11 N_CLKB_3 4.43756e-20
cc_305 N_MH_11 N_CLKB_29 0.000296768f
cc_306 N_MH_11 N_CLKB_24 0.000313017f
cc_307 N_MH_11 N_MM10_g 8.67603e-20
cc_308 N_MH_11 N_CLKB_23 0.000105619f
cc_309 N_MH_14 N_CLKB_23 0.00313943f
cc_310 N_MH_20 N_CLKB_24 0.000890644f
cc_311 N_MH_4 N_CLKB_2 0.000280209f
cc_312 N_MH_18 N_CLKB_25 0.000287173f
cc_313 N_MH_19 N_CLKB_23 0.000310499f
cc_314 N_MH_13 N_MM10_g 0.034246f
cc_315 N_MH_15 N_CLKB_24 0.000465454f
cc_316 N_MH_13 N_CLKB_2 0.000717753f
cc_317 N_MH_17 N_CLKB_24 0.000802909f
cc_318 N_MH_3 N_CLKB_1 0.000831729f
cc_319 N_MH_4 N_CLKB_24 0.000935401f
cc_320 N_MH_4 N_MM10_g 0.000955724f
cc_321 N_MH_3 N_MM4_g 0.0017231f
cc_322 N_MH_11 N_CLKB_1 0.00197805f
cc_323 N_MH_18 N_CLKB_29 0.00418313f
cc_324 N_MH_11 N_MM4_g 0.0347863f
cc_325 N_MH_1 N_MS_12 0.000875577f
cc_326 N_MM6_g N_MS_4 0.000917512f
cc_327 N_MH_18 N_MS_17 0.000959439f
cc_328 N_MH_1 N_MS_3 0.00263345f
cc_329 N_MM6_g N_MM11_g 0.00164916f
cc_330 N_MM6_g N_MS_5 0.00177411f
cc_331 N_MH_1 N_MS_14 0.00220504f
cc_332 N_MM6_g N_MS_14 0.0148237f
cc_333 N_MH_18 N_MS_16 0.00521426f
cc_334 N_MM6_g N_MS_12 0.0559548f
x_PM_SDFLx4_ASAP7_75t_R%PU1 VSS N_MM3_d N_MM2_d N_MM1_s N_PU1_8 N_PU1_2 N_PU1_7
+ N_PU1_1 N_PU1_9 PM_SDFLx4_ASAP7_75t_R%PU1
cc_335 N_PU1_8 N_CLKN_28 0.000180643f
cc_336 N_PU1_8 N_CLKN_2 0.000962632f
cc_337 N_PU1_2 N_MM1_g 0.000921045f
cc_338 N_PU1_8 N_MM1_g 0.0336828f
cc_339 N_PU1_7 N_SE_2 0.00065699f
cc_340 N_PU1_1 N_MM3_g 0.000914331f
cc_341 N_PU1_7 N_MM3_g 0.0338423f
cc_342 N_PU1_7 N_SI_1 0.000667145f
cc_343 N_PU1_1 N_MM2_g 0.000913388f
cc_344 N_PU1_7 N_MM2_g 0.0338386f
cc_345 N_PU1_9 N_CLKB_1 0.000405664f
cc_346 N_PU1_9 N_MM4_g 0.000495588f
cc_347 N_PU1_2 N_MM4_g 0.00047909f
cc_348 N_PU1_9 N_CLKB_29 0.000625553f
cc_349 N_PU1_9 N_CLKB_23 0.00154509f
cc_350 N_PU1_8 N_MH_13 0.00125228f
cc_351 N_PU1_2 N_MH_14 0.000661748f
cc_352 N_PU1_2 N_MH_19 0.000728006f
cc_353 N_PU1_9 N_MH_15 0.00112266f
cc_354 N_PU1_9 N_MH_19 0.00348599f
cc_355 N_PU1_2 N_MH_4 0.00462776f
cc_356 N_PU1_7 N_NET54_13 0.000560499f
cc_357 N_PU1_7 N_NET54_12 0.000640729f
cc_358 N_PU1_1 N_NET54_13 0.000664962f
cc_359 N_PU1_7 N_NET54_11 0.00112771f
cc_360 N_PU1_1 N_NET54_3 0.00185783f
cc_361 N_PU1_1 N_NET54_2 0.00429921f
cc_362 N_PU1_9 N_NET54_13 0.00959961f
x_PM_SDFLx4_ASAP7_75t_R%SI VSS SI N_MM2_g N_SI_9 N_SI_12 N_SI_8 N_SI_4 N_SI_1
+ N_SI_6 N_SI_5 N_SI_10 PM_SDFLx4_ASAP7_75t_R%SI
cc_363 N_SI_9 N_CLKN_23 9.01089e-20
cc_364 N_SI_12 N_CLKN_28 0.000269939f
cc_365 N_SI_8 N_CLKN_23 0.000999732f
cc_366 N_SI_9 N_CLKN_28 0.00318631f
cc_367 N_MM2_g N_SE_14 0.000233209f
cc_368 N_SI_4 N_SE_10 0.000608634f
cc_369 N_SI_1 N_SE_2 0.00210803f
cc_370 N_SI_9 N_SE_10 0.00111154f
cc_371 N_SI_9 N_SE_14 0.00151722f
cc_372 N_MM2_g N_MM3_g 0.00543449f
x_PM_SDFLx4_ASAP7_75t_R%NET54 VSS N_MM26_d N_MM0_d N_MM3_s N_MM2_s N_NET54_11
+ N_NET54_2 N_NET54_13 N_NET54_10 N_NET54_1 N_NET54_12 N_NET54_3
+ PM_SDFLx4_ASAP7_75t_R%NET54
cc_373 N_NET54_11 N_SE_2 0.00102735f
cc_374 N_NET54_2 N_MM3_g 0.000841639f
cc_375 N_NET54_13 N_SE_10 0.00240191f
cc_376 N_NET54_11 N_MM3_g 0.0335562f
cc_377 N_NET54_10 N_D_6 0.000725913f
cc_378 N_NET54_10 N_D_1 0.000786088f
cc_379 N_NET54_13 N_D_4 0.00135911f
cc_380 N_NET54_1 N_MM26_g 0.00185759f
cc_381 N_NET54_13 N_D_6 0.00227786f
cc_382 N_NET54_13 N_D_7 0.004737f
cc_383 N_NET54_10 N_MM26_g 0.034305f
cc_384 N_NET54_11 N_SEN_1 0.000924184f
cc_385 N_NET54_2 N_MM0_g 0.00086628f
cc_386 N_NET54_13 N_SEN_15 0.00224205f
cc_387 N_NET54_11 N_MM0_g 0.0344156f
cc_388 N_NET54_12 N_SI_1 0.000707847f
cc_389 N_NET54_3 N_MM2_g 0.000919355f
cc_390 N_NET54_13 N_SI_4 0.00214029f
cc_391 N_NET54_12 N_MM2_g 0.033747f
cc_392 N_NET54_12 N_CLKB_1 0.00100073f
cc_393 N_NET54_12 N_CLKB_23 0.000679536f
cc_394 N_NET54_3 N_MM4_g 0.0011783f
cc_395 N_NET54_13 N_CLKB_29 0.00391034f
cc_396 N_NET54_12 N_MM4_g 0.036224f
x_PM_SDFLx4_ASAP7_75t_R%SE VSS SE N_MM31_g N_MM3_g N_SE_15 N_SE_8 N_SE_12
+ N_SE_14 N_SE_10 N_SE_9 N_SE_7 N_SE_11 N_SE_1 N_SE_2 N_SE_13
+ PM_SDFLx4_ASAP7_75t_R%SE
cc_397 N_SE_15 N_CLKN_1 4.14287e-20
cc_398 N_SE_15 N_CLKN_22 6.37751e-20
cc_399 N_SE_8 N_CLKN_28 0.000163976f
cc_400 N_SE_12 N_CLKN_28 0.000175169f
cc_401 N_SE_14 N_CLKN_28 0.00019587f
cc_402 N_SE_10 N_CLKN_28 0.000835988f
cc_403 N_SE_9 N_CLKN_28 0.000326073f
cc_404 N_SE_7 N_CLKN_28 0.000814292f
cc_405 N_SE_15 N_CLKN_28 0.0287485f
x_PM_SDFLx4_ASAP7_75t_R%CLKN VSS N_MM23_g N_MM1_g N_MM12_g N_MM20_d N_MM21_d
+ N_CLKN_7 N_CLKN_26 N_CLKN_22 N_CLKN_1 N_CLKN_17 N_CLKN_21 N_CLKN_18 N_CLKN_19
+ N_CLKN_8 N_CLKN_28 N_CLKN_20 N_CLKN_16 N_CLKN_23 N_CLKN_2 N_CLKN_24 N_CLKN_3
+ N_CLKN_25 N_CLKN_27 PM_SDFLx4_ASAP7_75t_R%CLKN
cc_406 N_CLKN_7 N_MM20_g 0.00159706f
cc_407 N_CLKN_26 N_MM20_g 0.000248573f
cc_408 N_CLKN_22 N_MM20_g 0.000278047f
cc_409 N_CLKN_1 N_MM20_g 0.000381482f
cc_410 N_CLKN_17 N_MM20_g 0.0156456f
cc_411 N_CLKN_21 N_CLK_4 0.000462227f
cc_412 N_CLKN_18 N_CLK_5 0.000462891f
cc_413 N_CLKN_1 N_CLK_1 0.000473873f
cc_414 N_CLKN_19 N_CLK_4 0.000932105f
cc_415 N_CLKN_8 N_CLK_1 0.00115062f
cc_416 N_CLKN_28 N_CLK_5 0.00120808f
cc_417 N_CLKN_8 N_MM20_g 0.00137005f
cc_418 N_MM23_g N_MM20_g 0.00164693f
cc_419 N_CLKN_22 N_CLK_4 0.00200105f
cc_420 N_CLKN_17 N_CLK_1 0.00200609f
cc_421 N_CLKN_20 N_CLK_5 0.00394686f
cc_422 N_CLKN_26 N_CLK_4 0.00752557f
cc_423 N_CLKN_16 N_MM20_g 0.0555919f
x_PM_SDFLx4_ASAP7_75t_R%CLKB VSS N_MM4_g N_MM10_g N_MM13_g N_MM17_g N_MM22_d
+ N_MM23_d N_CLKB_10 N_CLKB_9 N_CLKB_29 N_CLKB_27 N_CLKB_22 N_CLKB_21 N_CLKB_1
+ N_CLKB_28 N_CLKB_26 N_CLKB_23 N_CLKB_4 N_CLKB_25 N_CLKB_20 N_CLKB_19
+ N_CLKB_24 N_CLKB_2 N_CLKB_3 PM_SDFLx4_ASAP7_75t_R%CLKB
cc_424 N_CLKB_10 N_CLK_5 0.000364571f
cc_425 N_CLKB_9 N_CLK_5 0.000147007f
cc_426 N_CLKB_29 N_CLK_5 5.55205e-20
cc_427 N_CLKB_27 N_CLK_5 8.13048e-20
cc_428 N_CLKB_22 N_CLK_5 0.000134975f
cc_429 N_CLKB_21 N_CLK_5 0.00121831f
cc_430 N_MM4_g N_CLKN_28 3.52501e-20
cc_431 N_CLKB_27 N_CLKN_19 6.05377e-20
cc_432 N_CLKB_1 N_CLKN_2 0.000142841f
cc_433 N_CLKB_9 N_MM23_g 0.00122293f
cc_434 N_CLKB_27 N_CLKN_21 8.10177e-20
cc_435 N_CLKB_28 N_CLKN_22 9.28534e-20
cc_436 N_CLKB_10 N_CLKN_22 0.000204781f
cc_437 N_CLKB_26 N_CLKN_24 0.00177607f
cc_438 N_CLKB_23 N_CLKN_28 0.000628452f
cc_439 N_CLKB_4 N_CLKN_3 0.000818871f
cc_440 N_CLKB_22 N_CLKN_22 0.00675599f
cc_441 N_CLKB_25 N_CLKN_28 0.000437184f
cc_442 N_CLKB_20 N_MM23_g 0.015767f
cc_443 N_CLKB_19 N_MM23_g 0.0537723f
cc_444 N_CLKB_29 N_CLKN_23 0.000527411f
cc_445 N_CLKB_24 N_CLKN_28 0.000549306f
cc_446 N_CLKB_27 N_CLKN_22 0.000603504f
cc_447 N_CLKB_2 N_CLKN_2 0.00159086f
cc_448 N_CLKB_10 N_CLKN_1 0.000749732f
cc_449 N_CLKB_22 N_CLKN_28 0.000813605f
cc_450 N_CLKB_29 N_CLKN_24 0.000883522f
cc_451 N_CLKB_21 N_CLKN_20 0.00096146f
cc_452 N_CLKB_3 N_CLKN_3 0.00237547f
cc_453 N_CLKB_10 N_MM23_g 0.00135834f
cc_454 N_MM17_g N_MM12_g 0.00163458f
cc_455 N_CLKB_20 N_CLKN_1 0.00172f
cc_456 N_MM10_g N_MM1_g 0.00335277f
cc_457 N_CLKB_24 N_CLKN_23 0.00425438f
cc_458 N_MM13_g N_MM12_g 0.00496365f
cc_459 N_CLKB_25 N_CLKN_24 0.00530411f
cc_460 N_CLKB_29 N_CLKN_28 0.073553f
cc_461 N_CLKB_10 N_SE_12 3.49832e-20
cc_462 N_CLKB_20 N_SE_12 4.67298e-20
cc_463 N_CLKB_19 N_SE_12 4.74871e-20
cc_464 N_MM4_g N_SE_12 5.13683e-20
cc_465 N_CLKB_21 N_SE_12 9.6634e-20
cc_466 N_CLKB_29 N_SE_12 0.000100729f
cc_467 N_CLKB_22 N_SE_1 0.000222109f
cc_468 N_CLKB_10 N_SE_8 0.000183594f
cc_469 N_CLKB_9 N_SE_7 0.000190076f
cc_470 N_CLKB_22 N_SE_8 0.00263121f
cc_471 N_CLKB_22 N_SE_7 0.00179416f
cc_472 N_CLKB_29 N_SE_9 0.000480469f
cc_473 N_CLKB_29 N_SE_10 0.00054126f
cc_474 N_CLKB_28 N_SE_11 0.00085695f
cc_475 N_CLKB_27 N_SE_13 0.000991394f
cc_476 N_CLKB_29 N_SE_15 0.00412702f
cc_477 N_CLKB_22 N_SE_12 0.00444164f
cc_478 N_CLKB_29 N_D_4 0.000746783f
cc_479 N_CLKB_29 N_D_7 0.00277794f
cc_480 N_CLKB_24 N_MM2_g 6.66654e-20
cc_481 N_CLKB_29 N_MM2_g 0.000173746f
cc_482 N_CLKB_23 N_MM2_g 0.000470375f
cc_483 N_CLKB_1 N_MM2_g 0.000207368f
cc_484 N_CLKB_23 N_SI_6 0.00026433f
cc_485 N_CLKB_23 N_SI_12 0.000300253f
cc_486 N_CLKB_1 N_SI_9 0.000310765f
cc_487 N_CLKB_1 N_SI_1 0.000966796f
cc_488 N_CLKB_29 N_SI_4 0.00132603f
cc_489 N_CLKB_23 N_SI_9 0.00175642f
cc_490 N_MM4_g N_MM2_g 0.00342403f
*END of SDFLx4_ASAP7_75t_R.pxi
.ENDS
** Design:	ASYNC_DFFHx1_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "ASYNC_DFFHx1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "ASYNC_DFFHx1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%NET077 VSS 2 4 1
c1 1 VSS 0.000858213f
r1 4 3 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9890 $Y=0.2160 $X2=0.9765 $Y2=0.2160
r2 2 1 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9550 $Y=0.2160 $X2=0.9595 $Y2=0.2160
r3 1 3 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9595 $Y=0.2160 $X2=0.9765 $Y2=0.2160
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.00861545f
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%PD1 VSS 2 4 1
c1 1 VSS 0.00100002f
r1 4 3 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3365 $Y2=0.0675
r2 2 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3195 $Y2=0.0675
r3 1 3 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3195 $Y=0.0675 $X2=0.3365 $Y2=0.0675
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.00945769f
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%CLK VSS 10 3 8 5 1 6 4 7
c1 1 VSS 0.00250274f
c2 3 VSS 0.0595942f
c3 4 VSS 0.00141499f
c4 5 VSS 0.00396291f
c5 6 VSS 0.00380145f
c6 7 VSS 0.00182501f
c7 8 VSS 0.00166788f
r1 6 20 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.2125 $X2=0.1080 $Y2=0.1910
r2 5 18 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0575 $X2=0.1080 $Y2=0.0790
r3 19 20 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.1910 $X2=0.1080 $Y2=0.1910
r4 8 16 2.66732 $w=1.57273e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1910 $X2=0.0810 $Y2=0.1745
r5 8 19 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1910 $X2=0.0945 $Y2=0.1910
r6 17 18 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.0790 $X2=0.1080 $Y2=0.0790
r7 7 13 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0790 $X2=0.0810 $Y2=0.0970
r8 7 17 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0790 $X2=0.0945 $Y2=0.0790
r9 15 16 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1645 $X2=0.0810 $Y2=0.1745
r10 14 15 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1530 $X2=0.0810 $Y2=0.1645
r11 12 14 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1530
r12 11 12 2.85657 $w=1.3e-08 $l=1.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1227 $X2=0.0810 $Y2=0.1350
r13 10 11 0.874462 $w=1.3e-08 $l=3.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1227
r14 10 4 1.57403 $w=1.3e-08 $l=6.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1122
r15 4 13 3.55614 $w=1.3e-08 $l=1.52e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1122 $X2=0.0810 $Y2=0.0970
r16 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r17 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%noxref_26 VSS 1
c1 1 VSS 0.0843809f
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%D VSS 21 3 6 4 1 5 8 9
c1 1 VSS 0.0102468f
c2 3 VSS 0.0830844f
c3 4 VSS 0.00399802f
c4 5 VSS 0.00350064f
c5 6 VSS 0.00174696f
c6 7 VSS 0.00733874f
c7 8 VSS 0.00110242f
c8 9 VSS 0.00723843f
r1 9 25 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2430 $Y2=0.2140
r2 7 23 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0360 $X2=0.2430 $Y2=0.0495
r3 24 25 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1850 $X2=0.2430 $Y2=0.2140
r4 5 8 3.60008 $w=1.51951e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.1555 $X2=0.2430 $Y2=0.1350
r5 5 24 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1555 $X2=0.2430 $Y2=0.1850
r6 21 22 2.2736 $w=1.3e-08 $l=9.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0820 $X2=0.2430 $Y2=0.0917
r7 21 20 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0820 $X2=0.2430 $Y2=0.0677
r8 20 23 4.25571 $w=1.3e-08 $l=1.82e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0677 $X2=0.2430 $Y2=0.0495
r9 19 22 4.25571 $w=1.3e-08 $l=1.83e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1100 $X2=0.2430 $Y2=0.0917
r10 18 19 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1195 $X2=0.2430 $Y2=0.1100
r11 4 8 1.61797 $w=1.675e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1230 $X2=0.2430 $Y2=0.1350
r12 4 18 0.816164 $w=1.3e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1230 $X2=0.2430 $Y2=0.1195
r13 16 17 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2715
+ $Y=0.1350 $X2=0.2810 $Y2=0.1350
r14 6 16 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2615
+ $Y=0.1350 $X2=0.2715 $Y2=0.1350
r15 6 8 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2615 $Y=0.1350 $X2=0.2430 $Y2=0.1350
r16 14 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2770 $Y=0.1350
+ $X2=0.2810 $Y2=0.1350
r17 12 14 4.43042 $w=1.53e-08 $l=7.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.2845 $Y=0.1350 $X2=0.2770 $Y2=0.1350
r18 1 11 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.2885
+ $Y=0.1350 $X2=0.2985 $Y2=0.1350
r19 1 12 1.86855 $w=1.78125e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.2885 $Y=0.1350 $X2=0.2845 $Y2=0.1350
r20 3 11 2.53453 $w=1.32811e-07 $l=1.5e-09 $layer=LIG $thickness=5.23243e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2985 $Y2=0.1350
r21 3 12 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2845 $Y2=0.1350
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%NET078 VSS 2 3 1
c1 1 VSS 0.000957754f
r1 2 1 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.2295 $X2=0.5940 $Y2=0.2295
r2 3 1 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.2295 $X2=0.5940 $Y2=0.2295
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%PD2 VSS 2 4 1
c1 1 VSS 0.000716587f
r1 4 3 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9350 $Y=0.2160 $X2=0.9305 $Y2=0.2160
r2 2 1 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9010 $Y=0.2160 $X2=0.9135 $Y2=0.2160
r3 1 3 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9135 $Y=0.2160 $X2=0.9305 $Y2=0.2160
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%NET076 VSS 2 3 1
c1 1 VSS 0.000859823f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0630 $Y=0.2160 $X2=1.0800 $Y2=0.2160
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0970 $Y=0.2160 $X2=1.0800 $Y2=0.2160
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%noxref_29 VSS 1
c1 1 VSS 0.0859164f
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%noxref_30 VSS 1
c1 1 VSS 0.0093487f
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%QN VSS 19 13 27 7 2 1 8 9
c1 1 VSS 0.00848947f
c2 2 VSS 0.00849608f
c3 7 VSS 0.0037691f
c4 8 VSS 0.00361315f
c5 9 VSS 0.00340801f
c6 10 VSS 0.00663835f
c7 11 VSS 0.00586406f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.3355 $Y=0.2025 $X2=1.3480 $Y2=0.2025
r2 27 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.3330 $Y=0.2025 $X2=1.3355 $Y2=0.2025
r3 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.3500 $Y=0.2025
+ $X2=1.3500 $Y2=0.2340
r4 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.3500
+ $Y=0.2340 $X2=1.3635 $Y2=0.2340
r5 11 22 7.56431 $w=1.42e-08 $l=3.75e-08 $layer=M1 $thickness=3.6e-08 $X=1.3770
+ $Y=0.2340 $X2=1.3770 $Y2=0.1965
r6 11 25 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3770 $Y=0.2340 $X2=1.3635 $Y2=0.2340
r7 21 22 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=1.3770
+ $Y=0.1675 $X2=1.3770 $Y2=0.1965
r8 20 21 2.04041 $w=1.3e-08 $l=8.8e-09 $layer=M1 $thickness=3.6e-08 $X=1.3770
+ $Y=0.1587 $X2=1.3770 $Y2=0.1675
r9 19 20 2.04041 $w=1.3e-08 $l=8.7e-09 $layer=M1 $thickness=3.6e-08 $X=1.3770
+ $Y=0.1500 $X2=1.3770 $Y2=0.1587
r10 19 18 7.05399 $w=1.3e-08 $l=3.03e-08 $layer=M1 $thickness=3.6e-08 $X=1.3770
+ $Y=0.1500 $X2=1.3770 $Y2=0.1197
r11 17 18 11.1348 $w=1.3e-08 $l=4.77e-08 $layer=M1 $thickness=3.6e-08 $X=1.3770
+ $Y=0.0720 $X2=1.3770 $Y2=0.1197
r12 9 16 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3770 $Y=0.0495 $X2=1.3770 $Y2=0.0360
r13 9 17 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.3770
+ $Y=0.0495 $X2=1.3770 $Y2=0.0720
r14 15 16 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.3635 $Y=0.0360 $X2=1.3770 $Y2=0.0360
r15 14 15 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.3500
+ $Y=0.0360 $X2=1.3635 $Y2=0.0360
r16 10 14 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.3385
+ $Y=0.0360 $X2=1.3500 $Y2=0.0360
r17 1 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.3500 $Y=0.0675
+ $X2=1.3500 $Y2=0.0360
r18 7 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.3355 $Y=0.0675 $X2=1.3480 $Y2=0.0675
r19 13 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.3330 $Y=0.0675 $X2=1.3355 $Y2=0.0675
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%SS VSS 13 14 30 44 45 3 15 4 7 9 1 16 6 8 5
c1 1 VSS 0.000217022f
c2 2 VSS 0.000757709f
c3 3 VSS 0.00237904f
c4 4 VSS 0.00606247f
c5 5 VSS 0.00167427f
c6 6 VSS 0.00136201f
c7 7 VSS 0.000341319f
c8 8 VSS 0.0045792f
c9 9 VSS 0.00111661f
c10 10 VSS 0.0014362f
c11 13 VSS 0.00599268f
c12 14 VSS 0.0220408f
c13 15 VSS 0.0035247f
c14 16 VSS 0.00306954f
r1 45 43 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.0970 $Y=0.0405 $X2=1.0945 $Y2=0.0405
r2 39 43 0.537037 $w=2.7e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.0800 $Y=0.0405 $X2=1.0945 $Y2=0.0405
r3 15 39 0.537037 $w=2.7e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.0655 $Y=0.0405 $X2=1.0800 $Y2=0.0405
r4 44 15 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.0630 $Y=0.0405 $X2=1.0655 $Y2=0.0405
r5 1 37 1.65643 $w=2.3e-08 $l=5e-09 $layer=LIG $thickness=4.8e-08 $X=0.9455
+ $Y=0.0910 $X2=0.9455 $Y2=0.0960
r6 13 1 1.9711 $w=1.43e-07 $l=4.40028e-08 $layer=LIG $thickness=5.27059e-08
+ $X=0.9450 $Y=0.1350 $X2=0.9455 $Y2=0.0910
r7 38 39 15.9139 $w=2.02e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.0800 $Y=0.0675 $X2=1.0800 $Y2=0.0405
r8 4 7 6.20751 $w=2.35778e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.0800 $Y=0.0825 $X2=1.0800 $Y2=0.0960
r9 4 38 8.84105 $w=2.02e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=1.0800
+ $Y=0.0825 $X2=1.0800 $Y2=0.0675
r10 36 37 14.7351 $w=2.02e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9590 $Y=0.0960 $X2=0.9455 $Y2=0.0960
r11 35 36 22.3973 $w=2.02e-08 $l=3.8e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9970 $Y=0.0960 $X2=0.9590 $Y2=0.0960
r12 34 35 8.84105 $w=2.02e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.0120 $Y=0.0960 $X2=0.9970 $Y2=0.0960
r13 33 34 8.25165 $w=2.02e-08 $l=1.4e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.0260 $Y=0.0960 $X2=1.0120 $Y2=0.0960
r14 32 33 8.25165 $w=2.02e-08 $l=1.4e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.0400 $Y=0.0960 $X2=1.0260 $Y2=0.0960
r15 31 32 7.95695 $w=2.02e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.0535 $Y=0.0960 $X2=1.0400 $Y2=0.0960
r16 3 7 6.20751 $w=2.35778e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.0665 $Y=0.0960 $X2=1.0800 $Y2=0.0960
r17 3 31 7.66224 $w=2.02e-08 $l=1.3e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.0665 $Y=0.0960 $X2=1.0535 $Y2=0.0960
r18 7 28 6.50222 $w=2.34571e-08 $l=1.4e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.0800 $Y=0.0960 $X2=1.0940 $Y2=0.0960
r19 16 25 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.1195 $Y=0.2160 $X2=1.1320 $Y2=0.2160
r20 30 16 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.1170 $Y=0.2160 $X2=1.1195 $Y2=0.2160
r21 27 28 7.95695 $w=2.02e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.1075 $Y=0.0960 $X2=1.0940 $Y2=0.0960
r22 26 27 7.66224 $w=2.02e-08 $l=1.3e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.1205 $Y=0.0960 $X2=1.1075 $Y2=0.0960
r23 5 9 9.60184 $w=2.6128e-08 $l=2.5e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.1340 $Y=0.0960 $X2=1.1590 $Y2=0.0960
r24 5 26 7.95695 $w=2.02e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.1340 $Y=0.0960 $X2=1.1205 $Y2=0.0960
r25 8 10 10.7315 $w=2.5e-08 $l=2.5e-08 $layer=LISD $thickness=2.7e-08 $X=1.1340
+ $Y=0.2010 $X2=1.1590 $Y2=0.2010
r26 8 25 14.1645 $w=2.18889e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.1340 $Y=0.2010 $X2=1.1340 $Y2=0.2280
r27 9 24 6.07417 $w=2.46e-08 $l=1.9e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.1590 $Y=0.0960 $X2=1.1590 $Y2=0.1150
r28 23 24 4.05162 $w=2.22e-08 $l=8e-09 $layer=LISD $thickness=2.7e-08 $X=1.1590
+ $Y=0.1230 $X2=1.1590 $Y2=0.1150
r29 22 23 6.07743 $w=2.22e-08 $l=1.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.1590 $Y=0.1350 $X2=1.1590 $Y2=0.1230
r30 21 22 5.82421 $w=2.22e-08 $l=1.15e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.1590 $Y=0.1465 $X2=1.1590 $Y2=0.1350
r31 20 21 4.05162 $w=2.22e-08 $l=8e-09 $layer=LISD $thickness=2.7e-08 $X=1.1590
+ $Y=0.1545 $X2=1.1590 $Y2=0.1465
r32 19 20 6.07743 $w=2.22e-08 $l=1.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.1590 $Y=0.1665 $X2=1.1590 $Y2=0.1545
r33 6 18 4.55807 $w=2.22e-08 $l=9.12414e-09 $layer=LISD $thickness=2.7e-08
+ $X=1.1590 $Y=0.1800 $X2=1.1605 $Y2=0.1890
r34 6 19 6.83711 $w=2.22e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.1590 $Y=0.1800 $X2=1.1590 $Y2=0.1665
r35 6 10 9.16613 $w=2.44455e-08 $l=2.1e-08 $layer=LISD $thickness=2.7e-08
+ $X=1.1590 $Y=0.1800 $X2=1.1590 $Y2=0.2010
r36 2 18 2.60296 $w=2.3e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08 $X=1.1605
+ $Y=0.2000 $X2=1.1605 $Y2=0.1890
r37 2 17 2.60296 $w=2.3e-08 $l=5e-10 $layer=LIG $thickness=4.8e-08 $X=1.1605
+ $Y=0.2000 $X2=1.1610 $Y2=0.2000
r38 2 10 8.01102 $w=2.45652e-08 $l=1.80278e-09 $layer=LISD
+ $thickness=3.70435e-08 $X=1.1605 $Y=0.2000 $X2=1.1590 $Y2=0.2010
r39 14 17 0.314665 $w=2.27e-07 $l=6.5e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.1610 $Y=0.1350 $X2=1.1610 $Y2=0.2000
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%noxref_28 VSS 1
c1 1 VSS 0.0090564f
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%SH VSS 12 13 69 71 76 80 14 5 23 15 18 17
+ 16 7 6 19 22 1 20 21 2
c1 1 VSS 0.000312365f
c2 2 VSS 0.00471478f
c3 5 VSS 0.00423007f
c4 6 VSS 0.00238243f
c5 7 VSS 0.00347981f
c6 12 VSS 0.0216525f
c7 13 VSS 0.0798918f
c8 14 VSS 0.00313136f
c9 15 VSS 0.00077759f
c10 16 VSS 0.00321222f
c11 17 VSS 0.00075956f
c12 18 VSS 0.00444996f
c13 19 VSS 0.00159349f
c14 20 VSS 0.00160122f
c15 21 VSS 0.00395933f
c16 22 VSS 0.00202943f
c17 23 VSS 0.0129237f
r1 80 79 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8810 $Y=0.0405 $X2=0.8785 $Y2=0.0405
r2 78 79 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8740 $Y=0.0405 $X2=0.8785 $Y2=0.0405
r3 5 78 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8620 $Y=0.0405 $X2=0.8740 $Y2=0.0405
r4 15 5 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.0405 $X2=0.8620 $Y2=0.0405
r5 14 5 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.0675 $X2=0.8620 $Y2=0.0675
r6 76 14 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.0675 $X2=0.8495 $Y2=0.0675
r7 5 65 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.0405
+ $X2=0.8670 $Y2=0.0390
r8 70 16 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8540 $Y=0.2295 $X2=0.8660 $Y2=0.2295
r9 17 70 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.2295 $X2=0.8540 $Y2=0.2295
r10 71 17 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.2295 $X2=0.8495 $Y2=0.2295
r11 69 68 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8810 $Y=0.2025 $X2=0.8785 $Y2=0.2025
r12 16 68 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8660 $Y=0.2025 $X2=0.8785 $Y2=0.2025
r13 65 66 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.8670
+ $Y=0.0390 $X2=0.8790 $Y2=0.0390
r14 64 66 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.0390 $X2=0.8790 $Y2=0.0390
r15 18 22 2.71097 $w=1.5e-08 $l=1.82483e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9090 $Y=0.0390 $X2=0.9270 $Y2=0.0420
r16 18 64 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.9090
+ $Y=0.0390 $X2=0.8910 $Y2=0.0390
r17 7 16 14.1645 $w=2.18889e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8640 $Y=0.2010 $X2=0.8640 $Y2=0.2280
r18 2 55 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.3230 $Y=0.1350
+ $X2=1.3230 $Y2=0.1440
r19 13 2 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=1.3230
+ $Y=0.1350 $X2=1.3230 $Y2=0.1350
r20 22 51 1.31184 $w=1.63333e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.9270 $Y=0.0420 $X2=0.9270 $Y2=0.0510
r21 6 58 17.6821 $w=2.02e-08 $l=3e-08 $layer=LISD $thickness=2.7e-08 $X=0.8970
+ $Y=0.2010 $X2=0.9270 $Y2=0.2010
r22 6 7 17.7009 $w=2.15818e-08 $l=3.3e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8970 $Y=0.2010 $X2=0.8640 $Y2=0.2010
r23 21 55 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=1.3230
+ $Y=0.1145 $X2=1.3230 $Y2=0.1440
r24 50 51 1.16595 $w=1.3e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.9270
+ $Y=0.0560 $X2=0.9270 $Y2=0.0510
r25 49 50 1.51573 $w=1.3e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.9270
+ $Y=0.0625 $X2=0.9270 $Y2=0.0560
r26 48 49 1.63233 $w=1.3e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.9270
+ $Y=0.0695 $X2=0.9270 $Y2=0.0625
r27 47 48 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.9270
+ $Y=0.0810 $X2=0.9270 $Y2=0.0695
r28 46 47 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.9270
+ $Y=0.0935 $X2=0.9270 $Y2=0.0810
r29 45 58 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.9270 $Y=0.1975
+ $X2=0.9270 $Y2=0.2010
r30 44 45 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.9270
+ $Y=0.1770 $X2=0.9270 $Y2=0.1975
r31 43 44 5.59655 $w=1.3e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.9270
+ $Y=0.1530 $X2=0.9270 $Y2=0.1770
r32 19 43 7.57867 $w=1.3e-08 $l=3.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.9270
+ $Y=0.1205 $X2=0.9270 $Y2=0.1530
r33 19 46 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9270
+ $Y=0.1205 $X2=0.9270 $Y2=0.0935
r34 41 55 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=1.3230 $Y=0.1530
+ $X2=1.3230 $Y2=0.1440
r35 40 41 15.6237 $w=1.3e-08 $l=6.7e-08 $layer=M2 $thickness=3.6e-08 $X=1.2560
+ $Y=0.1530 $X2=1.3230 $Y2=0.1530
r36 39 40 23.0858 $w=1.3e-08 $l=9.9e-08 $layer=M2 $thickness=3.6e-08 $X=1.1570
+ $Y=0.1530 $X2=1.2560 $Y2=0.1530
r37 38 39 11.6595 $w=1.3e-08 $l=5e-08 $layer=M2 $thickness=3.6e-08 $X=1.1070
+ $Y=0.1530 $X2=1.1570 $Y2=0.1530
r38 37 38 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=1.0825
+ $Y=0.1530 $X2=1.1070 $Y2=0.1530
r39 33 34 9.56078 $w=1.3e-08 $l=4.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.9310
+ $Y=0.1530 $X2=0.9720 $Y2=0.1530
r40 33 43 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.9310 $Y=0.1530
+ $X2=0.9270 $Y2=0.1530
r41 23 34 15.2739 $w=1.3e-08 $l=6.55e-08 $layer=M2 $thickness=3.6e-08 $X=1.0375
+ $Y=0.1530 $X2=0.9720 $Y2=0.1530
r42 23 37 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M2 $thickness=3.6e-08 $X=1.0375
+ $Y=0.1530 $X2=1.0825 $Y2=0.1530
r43 30 38 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=1.1070 $Y=0.1440
+ $X2=1.1070 $Y2=0.1530
r44 20 30 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=1.1070
+ $Y=0.1145 $X2=1.1070 $Y2=0.1440
r45 12 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=1.1070
+ $Y=0.1350 $X2=1.1070 $Y2=0.1350
r46 1 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.1070 $Y=0.1350
+ $X2=1.1070 $Y2=0.1440
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%NET079 VSS 2 3 1
c1 1 VSS 0.000829673f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.2160 $X2=0.7020 $Y2=0.2160
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.2160 $X2=0.7020 $Y2=0.2160
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%NET051 VSS 7 11 4 5 1
c1 1 VSS 0.00700205f
c2 4 VSS 0.00189002f
c3 5 VSS 0.00224118f
r1 11 10 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.2295 $X2=0.5545 $Y2=0.2295
r2 5 10 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5420 $Y=0.2295 $X2=0.5545 $Y2=0.2295
r3 8 5 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08 $X=0.5130
+ $Y=0.2295 $X2=0.5400 $Y2=0.2295
r4 1 8 12.6992 $w=2.32e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08 $X=0.4860
+ $Y=0.2295 $X2=0.5130 $Y2=0.2295
r5 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2295 $X2=0.4840 $Y2=0.2295
r6 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2295 $X2=0.4715 $Y2=0.2295
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%RESET VSS 24 5 6 12 10 7 8 2 9 11 1
c1 1 VSS 0.00321126f
c2 2 VSS 0.00179614f
c3 5 VSS 0.0608868f
c4 6 VSS 0.0496184f
c5 7 VSS 0.00077689f
c6 8 VSS 0.00124738f
c7 9 VSS 0.00226846f
c8 10 VSS 0.00203018f
c9 11 VSS 0.000769163f
c10 12 VSS 0.00151691f
r1 8 11 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.6460
+ $Y=0.1890 $X2=0.6210 $Y2=0.1890
r2 11 35 1.84873 $w=1.888e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1890 $X2=0.6210 $Y2=0.1740
r3 1 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6210 $Y=0.1590
+ $X2=0.6210 $Y2=0.1570
r4 5 1 2.92627 $w=1.245e-07 $l=2.4e-08 $layer=LIG $thickness=5.2e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1590
r5 34 35 1.86552 $w=1.3e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1660 $X2=0.6210 $Y2=0.1740
r6 33 34 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1570 $X2=0.6210 $Y2=0.1660
r7 7 33 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1380 $X2=0.6210 $Y2=0.1570
r8 7 32 3.71668 $w=1.51429e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.1380 $X2=0.6210 $Y2=0.1170
r9 10 30 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6335
+ $Y=0.1170 $X2=0.6460 $Y2=0.1170
r10 10 32 1.73456 $w=1.66e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6335 $Y=0.1170 $X2=0.6210 $Y2=0.1170
r11 28 29 13.4084 $w=1.3e-08 $l=5.75e-08 $layer=M2 $thickness=3.6e-08 $X=0.6460
+ $Y=0.1170 $X2=0.7035 $Y2=0.1170
r12 28 30 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.6460 $Y=0.1170
+ $X2=0.6460 $Y2=0.1170
r13 26 29 14.9241 $w=1.3e-08 $l=6.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.7675
+ $Y=0.1170 $X2=0.7035 $Y2=0.1170
r14 24 25 2.85657 $w=1.3e-08 $l=1.22e-08 $layer=M2 $thickness=3.6e-08 $X=0.8280
+ $Y=0.1170 $X2=0.8402 $Y2=0.1170
r15 24 23 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M2 $thickness=3.6e-08 $X=0.8280
+ $Y=0.1170 $X2=0.8052 $Y2=0.1170
r16 23 26 8.80291 $w=1.3e-08 $l=3.77e-08 $layer=M2 $thickness=3.6e-08 $X=0.8052
+ $Y=0.1170 $X2=0.7675 $Y2=0.1170
r17 22 25 9.85227 $w=1.3e-08 $l=4.23e-08 $layer=M2 $thickness=3.6e-08 $X=0.8825
+ $Y=0.1170 $X2=0.8402 $Y2=0.1170
r18 12 20 17.3726 $w=1.3e-08 $l=7.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.9785
+ $Y=0.1170 $X2=1.0530 $Y2=0.1170
r19 12 22 22.3862 $w=1.3e-08 $l=9.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.9785
+ $Y=0.1170 $X2=0.8825 $Y2=0.1170
r20 18 20 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=1.0530 $Y=0.1260
+ $X2=1.0530 $Y2=0.1170
r21 9 18 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1055 $X2=1.0530 $Y2=0.1260
r22 6 2 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=1.0530
+ $Y=0.1350 $X2=1.0530 $Y2=0.1350
r23 2 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=1.0530 $Y=0.1350
+ $X2=1.0530 $Y2=0.1260
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%PU1 VSS 7 10 5 4 1
c1 1 VSS 0.0102147f
c2 4 VSS 0.00317726f
c3 5 VSS 0.00183678f
r1 10 9 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r2 8 9 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r3 5 8 0.123457 $w=8.1e-08 $l=1e-08 $layer=P_src_drn $thickness=1e-09 $X=0.3780
+ $Y=0.2025 $X2=0.3880 $Y2=0.2025
r4 4 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3220 $Y2=0.2025
r5 7 4 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r6 1 5 1e-05
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%NET020 VSS 11 25 26 7 1 8 2 9
c1 1 VSS 0.00498693f
c2 2 VSS 0.00925891f
c3 7 VSS 0.0022953f
c4 8 VSS 0.00430531f
c5 9 VSS 0.0199439f
r1 26 24 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.0540 $X2=0.6085 $Y2=0.0540
r2 2 24 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.0540 $X2=0.6085 $Y2=0.0540
r3 8 2 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.0540 $X2=0.5940 $Y2=0.0540
r4 25 8 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0540 $X2=0.5795 $Y2=0.0540
r5 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0540
+ $X2=0.5940 $Y2=0.0360
r6 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5805
+ $Y=0.0360 $X2=0.5940 $Y2=0.0360
r7 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0360 $X2=0.5805 $Y2=0.0360
r8 18 19 3.38125 $w=1.3e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.5525
+ $Y=0.0360 $X2=0.5670 $Y2=0.0360
r9 17 18 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.5165
+ $Y=0.0360 $X2=0.5525 $Y2=0.0360
r10 16 17 9.211 $w=1.3e-08 $l=3.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4770
+ $Y=0.0360 $X2=0.5165 $Y2=0.0360
r11 15 16 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0360 $X2=0.4770 $Y2=0.0360
r12 14 15 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4455
+ $Y=0.0360 $X2=0.4590 $Y2=0.0360
r13 13 14 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4455 $Y2=0.0360
r14 12 13 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4205
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r15 9 12 0.932759 $w=1.3e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.4165
+ $Y=0.0360 $X2=0.4205 $Y2=0.0360
r16 1 13 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0540
+ $X2=0.4320 $Y2=0.0360
r17 7 1 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0540 $X2=0.4300 $Y2=0.0540
r18 11 7 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0540 $X2=0.4175 $Y2=0.0540
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%noxref_27 VSS 1
c1 1 VSS 0.0357567f
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%CLKN VSS 15 16 17 18 90 92 28 10 9 20 19 1
+ 23 22 27 29 21 30 24 2 25 26 4 3
c1 1 VSS 0.00186252f
c2 2 VSS 0.000397928f
c3 3 VSS 0.000313519f
c4 4 VSS 0.000175258f
c5 9 VSS 0.00787276f
c6 10 VSS 0.00791152f
c7 15 VSS 0.0591836f
c8 16 VSS 0.00535461f
c9 17 VSS 0.00554667f
c10 18 VSS 0.004532f
c11 19 VSS 0.00705163f
c12 20 VSS 0.00697718f
c13 21 VSS 0.00637697f
c14 22 VSS 0.00406351f
c15 23 VSS 0.000796715f
c16 24 VSS 0.000680733f
c17 25 VSS 0.000187943f
c18 26 VSS 0.000334127f
c19 27 VSS 0.00761169f
c20 28 VSS 0.00183687f
c21 29 VSS 0.00686874f
c22 30 VSS 0.0224712f
r1 92 91 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r2 20 91 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r3 90 89 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r4 19 89 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r5 10 86 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0550 $Y2=0.2340
r6 9 82 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0550 $Y2=0.0360
r7 15 76 0.314665 $w=2.27e-07 $l=0 $layer=Gate_1 $thickness=5.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r8 85 86 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.2340 $X2=0.0550 $Y2=0.2340
r9 84 85 1.28254 $w=1.3e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.2340 $X2=0.0460 $Y2=0.2340
r10 29 72 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0270 $Y2=0.2125
r11 29 84 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0405 $Y2=0.2340
r12 81 82 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.0360 $X2=0.0550 $Y2=0.0360
r13 80 81 1.28254 $w=1.3e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.0360 $X2=0.0460 $Y2=0.0360
r14 27 70 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0360 $X2=0.0270 $Y2=0.0575
r15 27 80 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0360 $X2=0.0405 $Y2=0.0360
r16 74 75 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.1335
+ $Y=0.1350 $X2=0.1435 $Y2=0.1350
r17 74 76 2.21986 $w=2.2e-08 $l=1.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1335
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r18 1 75 1.86855 $w=1.78125e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1475 $Y=0.1350 $X2=0.1435 $Y2=0.1350
r19 1 78 4.43042 $w=1.53e-08 $l=7.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1475
+ $Y=0.1350 $X2=0.1550 $Y2=0.1350
r20 71 72 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1910 $X2=0.0270 $Y2=0.2125
r21 22 28 2.9164 $w=1.82105e-08 $l=1.978e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1720 $X2=0.0325 $Y2=0.1530
r22 22 71 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1720 $X2=0.0270 $Y2=0.1910
r23 69 70 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0790 $X2=0.0270 $Y2=0.0575
r24 21 28 7.11381 $w=1.56757e-08 $l=3.74066e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1160 $X2=0.0325 $Y2=0.1530
r25 21 69 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1160 $X2=0.0270 $Y2=0.0790
r26 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
r27 16 2 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r28 3 57 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1350
+ $X2=0.4590 $Y2=0.1440
r29 17 3 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r30 63 78 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1510 $Y=0.1440
+ $X2=0.1550 $Y2=0.1350
r31 23 63 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1510
+ $Y=0.1160 $X2=0.1510 $Y2=0.1440
r32 28 53 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.0325 $Y=0.1530
+ $X2=0.0330 $Y2=0.1530
r33 24 61 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1530
r34 25 57 4.89699 $w=1.3e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1230 $X2=0.4590 $Y2=0.1440
r35 55 56 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M2 $thickness=3.6e-08 $X=0.1510
+ $Y=0.1530 $X2=0.1675 $Y2=0.1530
r36 55 63 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1510 $Y=0.1530
+ $X2=0.1510 $Y2=0.1440
r37 54 55 13.7582 $w=1.3e-08 $l=5.9e-08 $layer=M2 $thickness=3.6e-08 $X=0.0920
+ $Y=0.1530 $X2=0.1510 $Y2=0.1530
r38 53 54 13.7582 $w=1.3e-08 $l=5.9e-08 $layer=M2 $thickness=3.6e-08 $X=0.0330
+ $Y=0.1530 $X2=0.0920 $Y2=0.1530
r39 50 51 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1530 $X2=0.3620 $Y2=0.1530
r40 50 61 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.3510 $Y=0.1530
+ $X2=0.3510 $Y2=0.1530
r41 49 50 21.5701 $w=1.3e-08 $l=9.25e-08 $layer=M2 $thickness=3.6e-08 $X=0.2585
+ $Y=0.1530 $X2=0.3510 $Y2=0.1530
r42 49 56 21.2203 $w=1.3e-08 $l=9.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.2585
+ $Y=0.1530 $X2=0.1675 $Y2=0.1530
r43 47 48 21.2203 $w=1.3e-08 $l=9.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1530 $X2=0.5500 $Y2=0.1530
r44 47 57 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4590 $Y=0.1530
+ $X2=0.4590 $Y2=0.1440
r45 46 47 12.1259 $w=1.3e-08 $l=5.2e-08 $layer=M2 $thickness=3.6e-08 $X=0.4070
+ $Y=0.1530 $X2=0.4590 $Y2=0.1530
r46 46 51 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M2 $thickness=3.6e-08 $X=0.4070
+ $Y=0.1530 $X2=0.3620 $Y2=0.1530
r47 30 44 25.0679 $w=1.3e-08 $l=1.075e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.7305 $Y=0.1530 $X2=0.8380 $Y2=0.1530
r48 30 48 42.0908 $w=1.3e-08 $l=1.805e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.7305 $Y=0.1530 $X2=0.5500 $Y2=0.1530
r49 42 44 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.8380 $Y=0.1530
+ $X2=0.8380 $Y2=0.1530
r50 41 42 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.8380
+ $Y=0.1330 $X2=0.8380 $Y2=0.1530
r51 40 41 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.8380
+ $Y=0.1130 $X2=0.8380 $Y2=0.1330
r52 26 40 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.8380
+ $Y=0.1015 $X2=0.8380 $Y2=0.1130
r53 4 37 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.8370
+ $Y=0.1110 $X2=0.8370 $Y2=0.1110
r54 4 40 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8370 $Y=0.1110
+ $X2=0.8380 $Y2=0.1130
r55 18 37 0.314665 $w=2.27e-07 $l=2.4e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.8370 $Y=0.1350 $X2=0.8370 $Y2=0.1110
r56 10 20 1e-05
r57 9 19 1e-05
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%PD3 VSS 15 18 29 7 1 11 9 10 8 2
c1 1 VSS 0.00576357f
c2 2 VSS 0.00572267f
c3 7 VSS 0.00330097f
c4 8 VSS 0.00323752f
c5 9 VSS 0.00437594f
c6 10 VSS 0.00458857f
c7 11 VSS 0.0118224f
r1 8 2 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.1735 $Y=0.0405 $X2=1.1860 $Y2=0.0405
r2 29 8 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.1710 $Y=0.0405 $X2=1.1735 $Y2=0.0405
r3 2 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.1880 $Y=0.0405
+ $X2=1.1860 $Y2=0.0450
r4 10 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.1725
+ $Y=0.0450 $X2=1.1860 $Y2=0.0450
r5 24 26 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=1.1840 $Y=0.0450 $X2=1.1860
+ $Y2=0.0450
r6 23 24 14.691 $w=1.3e-08 $l=6.3e-08 $layer=M2 $thickness=3.6e-08 $X=1.1210
+ $Y=0.0450 $X2=1.1840 $Y2=0.0450
r7 22 23 43.0235 $w=1.3e-08 $l=1.845e-07 $layer=M2 $thickness=3.6e-08 $X=0.9365
+ $Y=0.0450 $X2=1.1210 $Y2=0.0450
r8 21 22 32.53 $w=1.3e-08 $l=1.395e-07 $layer=M2 $thickness=3.6e-08 $X=0.7970
+ $Y=0.0450 $X2=0.9365 $Y2=0.0450
r9 11 21 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.7855
+ $Y=0.0450 $X2=0.7970 $Y2=0.0450
r10 19 21 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.7995 $Y=0.0450
+ $X2=0.7970 $Y2=0.0450
r11 9 19 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.0450 $X2=0.7995 $Y2=0.0450
r12 1 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8100 $Y=0.0540
+ $X2=0.7995 $Y2=0.0450
r13 18 17 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8270 $Y=0.0540 $X2=0.8245 $Y2=0.0540
r14 1 17 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8120 $Y=0.0540 $X2=0.8245 $Y2=0.0540
r15 14 1 0.222222 $w=5.4e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8000 $Y=0.0540 $X2=0.8120 $Y2=0.0540
r16 7 14 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.0540 $X2=0.8000 $Y2=0.0540
r17 15 7 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.0540 $X2=0.7955 $Y2=0.0540
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%MH VSS 9 53 54 76 80 13 18 1 11 15 14 10 19
+ 16 20 3 17 4 22 21
c1 1 VSS 0.0032375f
c2 3 VSS 0.00476806f
c3 4 VSS 0.00493941f
c4 9 VSS 0.0321873f
c5 10 VSS 0.00247756f
c6 11 VSS 0.000620847f
c7 12 VSS 6.1547e-20
c8 13 VSS 0.00215879f
c9 14 VSS 8.90325e-20
c10 15 VSS 0.00243637f
c11 16 VSS 0.00587139f
c12 17 VSS 0.000991312f
c13 18 VSS 0.00124044f
c14 19 VSS 0.0013751f
c15 20 VSS 0.000295687f
c16 21 VSS 0.00225081f
c17 22 VSS 0.00635594f
r1 80 79 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2295 $X2=0.4465 $Y2=0.2295
r2 78 79 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4420 $Y=0.2295 $X2=0.4465 $Y2=0.2295
r3 4 78 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4300 $Y=0.2295 $X2=0.4420 $Y2=0.2295
r4 14 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2295 $X2=0.4300 $Y2=0.2295
r5 13 4 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.1890 $X2=0.4300 $Y2=0.1890
r6 76 13 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.1890 $X2=0.4175 $Y2=0.1890
r7 4 70 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2295
+ $X2=0.4320 $Y2=0.2340
r8 70 71 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4455 $Y2=0.2340
r9 68 71 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4455 $Y2=0.2340
r10 16 21 2.55791 $w=1.46667e-08 $l=1.8554e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4770 $Y=0.2340 $X2=0.4950 $Y2=0.2295
r11 16 68 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4770
+ $Y=0.2340 $X2=0.4590 $Y2=0.2340
r12 21 66 3.02429 $w=1.44516e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4950 $Y=0.2295 $X2=0.4950 $Y2=0.2140
r13 65 66 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4950
+ $Y=0.1850 $X2=0.4950 $Y2=0.2140
r14 64 65 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4950
+ $Y=0.1655 $X2=0.4950 $Y2=0.1850
r15 63 64 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4950
+ $Y=0.1450 $X2=0.4950 $Y2=0.1655
r16 62 63 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4950
+ $Y=0.1225 $X2=0.4950 $Y2=0.1450
r17 61 62 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4950
+ $Y=0.1135 $X2=0.4950 $Y2=0.1225
r18 60 61 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4950
+ $Y=0.1045 $X2=0.4950 $Y2=0.1135
r19 17 20 1.73214 $w=1.90828e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4950 $Y=0.0955 $X2=0.4950 $Y2=0.0810
r20 17 60 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4950
+ $Y=0.0955 $X2=0.4950 $Y2=0.1045
r21 58 59 0.264706 $w=1.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.0725 $X2=0.3925 $Y2=0.0725
r22 11 58 0.705882 $w=1.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3760 $Y=0.0725 $X2=0.3880 $Y2=0.0725
r23 12 11 0.735294 $w=1.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.0725 $X2=0.3760 $Y2=0.0725
r24 54 52 0.0675676 $w=3.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0455 $X2=0.3925 $Y2=0.0455
r25 11 52 0.391892 $w=3.7e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.0455 $X2=0.3925 $Y2=0.0455
r26 11 59 0.471383 $w=3.35517e-08 $l=3.06472e-08 $layer=N_src_drn
+ $thickness=1e-09 $X=0.3780 $Y=0.0455 $X2=0.3925 $Y2=0.0725
r27 10 11 0.391892 $w=3.7e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.0455 $X2=0.3780 $Y2=0.0455
r28 53 10 0.0675676 $w=3.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0455 $X2=0.3635 $Y2=0.0455
r29 3 11 16.798 $w=2.02e-08 $l=2.85e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.3780 $Y=0.0825 $X2=0.3780 $Y2=0.0540
r30 3 49 5.59933 $w=2.02e-08 $l=9.5e-09 $layer=LISD $thickness=2.7e-08
+ $X=0.3780 $Y=0.0825 $X2=0.3780 $Y2=0.0920
r31 18 46 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5080
+ $Y=0.0810 $X2=0.5210 $Y2=0.0810
r32 18 20 1.38235 $w=1.64615e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5080 $Y=0.0810 $X2=0.4950 $Y2=0.0810
r33 44 49 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.0830
+ $X2=0.3780 $Y2=0.0920
r34 15 44 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0630 $X2=0.3780 $Y2=0.0830
r35 42 43 13.9914 $w=1.3e-08 $l=6e-08 $layer=M2 $thickness=3.6e-08 $X=0.5210
+ $Y=0.0810 $X2=0.5810 $Y2=0.0810
r36 42 46 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.5210 $Y=0.0810
+ $X2=0.5210 $Y2=0.0810
r37 41 42 16.6731 $w=1.3e-08 $l=7.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.4495
+ $Y=0.0810 $X2=0.5210 $Y2=0.0810
r38 40 41 16.6731 $w=1.3e-08 $l=7.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0810 $X2=0.4495 $Y2=0.0810
r39 40 44 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.3780 $Y=0.0810
+ $X2=0.3780 $Y2=0.0830
r40 22 37 13.4084 $w=1.3e-08 $l=5.75e-08 $layer=M2 $thickness=3.6e-08 $X=0.6805
+ $Y=0.0810 $X2=0.7380 $Y2=0.0810
r41 22 43 23.2024 $w=1.3e-08 $l=9.95e-08 $layer=M2 $thickness=3.6e-08 $X=0.6805
+ $Y=0.0810 $X2=0.5810 $Y2=0.0810
r42 34 35 3.38125 $w=1.3e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.7380
+ $Y=0.0955 $X2=0.7380 $Y2=0.1100
r43 19 34 3.38125 $w=1.3e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.7380
+ $Y=0.0810 $X2=0.7380 $Y2=0.0955
r44 19 37 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.7380 $Y=0.0810
+ $X2=0.7380 $Y2=0.0810
r45 28 30 2.1068 $w=2.17667e-08 $l=7.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.7340 $Y=0.1100 $X2=0.7415 $Y2=0.1100
r46 28 35 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7340 $Y=0.1100
+ $X2=0.7380 $Y2=0.1100
r47 1 28 2.1415 $w=2.4e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.7240
+ $Y=0.1100 $X2=0.7340 $Y2=0.1100
r48 1 29 1.27796 $w=2.33909e-08 $l=5.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.7240 $Y=0.1100 $X2=0.7185 $Y2=0.1100
r49 27 28 1.07075 $w=2.4e-08 $l=5e-09 $layer=LIG $thickness=4.8e-08 $X=0.7290
+ $Y=0.1100 $X2=0.7340 $Y2=0.1100
r50 27 29 0.207209 $w=1.73e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7290 $Y=0.1100 $X2=0.7185 $Y2=0.1100
r51 27 30 1.03605 $w=1.73e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7290 $Y=0.1100 $X2=0.7415 $Y2=0.1100
r52 9 27 0.314665 $w=2.27e-07 $l=2.5e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.7290 $Y=0.1350 $X2=0.7290 $Y2=0.1100
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%SET VSS 51 7 8 9 12 11 5 10 1 3
c1 1 VSS 0.00118098f
c2 2 VSS 0.00121099f
c3 3 VSS 0.00126572f
c4 5 VSS 0.00552469f
c5 7 VSS 0.0607486f
c6 8 VSS 0.0320003f
c7 9 VSS 0.0493664f
c8 10 VSS 0.00106155f
c9 11 VSS 0.00182333f
c10 12 VSS 0.00172783f
r1 51 50 4.37231 $w=1.3e-08 $l=1.88e-08 $layer=M2 $thickness=3.6e-08 $X=0.8430
+ $Y=0.0810 $X2=0.8242 $Y2=0.0810
r2 49 50 6.35442 $w=1.3e-08 $l=2.72e-08 $layer=M2 $thickness=3.6e-08 $X=0.7970
+ $Y=0.0810 $X2=0.8242 $Y2=0.0810
r3 12 49 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.7855
+ $Y=0.0810 $X2=0.7970 $Y2=0.0810
r4 46 49 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.7990 $Y=0.0810 $X2=0.7970
+ $Y2=0.0810
r5 45 46 1.83642 $w=1.41111e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.7900
+ $Y=0.0810 $X2=0.7990 $Y2=0.0810
r6 44 45 0.714311 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.0810 $X2=0.7900 $Y2=0.0810
r7 11 39 1.02025 $w=1.48182e-08 $l=1.43265e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7760 $Y=0.0810 $X2=0.7830 $Y2=0.0935
r8 11 44 0.714311 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.7760
+ $Y=0.0810 $X2=0.7830 $Y2=0.0810
r9 1 35 2.60296 $w=2.3e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.6755
+ $Y=0.1590 $X2=0.6755 $Y2=0.1590
r10 7 1 2.91763 $w=1.20143e-07 $l=2.40052e-08 $layer=LIG $thickness=5.18095e-08
+ $X=0.6750 $Y=0.1350 $X2=0.6755 $Y2=0.1590
r11 38 39 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.0980 $X2=0.7830 $Y2=0.0935
r12 37 38 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1160 $X2=0.7830 $Y2=0.0980
r13 10 36 3.96423 $w=1.3e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1415 $X2=0.7830 $Y2=0.1585
r14 10 37 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1415 $X2=0.7830 $Y2=0.1160
r15 2 27 8.43855 $w=2.12286e-08 $l=0 $layer=LISD $thickness=3.9e-08 $X=0.7830
+ $Y=0.1590 $X2=0.7830 $Y2=0.1590
r16 2 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7830 $Y=0.1590
+ $X2=0.7830 $Y2=0.1585
r17 8 2 3.44859 $w=1.15182e-07 $l=2.4e-08 $layer=LIG $thickness=5.16364e-08
+ $X=0.7830 $Y=0.1350 $X2=0.7830 $Y2=0.1590
r18 34 35 7.66224 $w=2.02e-08 $l=1.5e-09 $layer=LISD $thickness=2.7e-08
+ $X=0.6770 $Y=0.1590 $X2=0.6755 $Y2=0.1590
r19 33 34 14.7351 $w=2.02e-08 $l=2.5e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7020 $Y=0.1590 $X2=0.6770 $Y2=0.1590
r20 32 33 8.25165 $w=2.02e-08 $l=1.4e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7160 $Y=0.1590 $X2=0.7020 $Y2=0.1590
r21 31 32 8.84105 $w=2.02e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7310 $Y=0.1590 $X2=0.7160 $Y2=0.1590
r22 30 31 10.904 $w=2.02e-08 $l=1.85e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7495 $Y=0.1590 $X2=0.7310 $Y2=0.1590
r23 29 30 7.07284 $w=2.02e-08 $l=1.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7615 $Y=0.1590 $X2=0.7495 $Y2=0.1590
r24 27 28 7.07284 $w=2.02e-08 $l=1.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7830 $Y=0.1590 $X2=0.7950 $Y2=0.1590
r25 27 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7830 $Y=0.1590
+ $X2=0.7830 $Y2=0.1585
r26 26 27 7.07284 $w=2.02e-08 $l=1.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7710 $Y=0.1590 $X2=0.7830 $Y2=0.1590
r27 26 29 5.59933 $w=2.02e-08 $l=9.5e-09 $layer=LISD $thickness=2.7e-08
+ $X=0.7710 $Y=0.1590 $X2=0.7615 $Y2=0.1590
r28 25 28 8.84105 $w=2.02e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8100 $Y=0.1590 $X2=0.7950 $Y2=0.1590
r29 24 25 8.25165 $w=2.02e-08 $l=1.4e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8240 $Y=0.1590 $X2=0.8100 $Y2=0.1590
r30 23 24 7.95695 $w=2.02e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8375 $Y=0.1590 $X2=0.8240 $Y2=0.1590
r31 22 23 7.66224 $w=2.02e-08 $l=1.3e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8505 $Y=0.1590 $X2=0.8375 $Y2=0.1590
r32 21 22 7.95695 $w=2.02e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8640 $Y=0.1590 $X2=0.8505 $Y2=0.1590
r33 20 21 8.25165 $w=2.02e-08 $l=1.4e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8780 $Y=0.1590 $X2=0.8640 $Y2=0.1590
r34 19 20 7.95695 $w=2.02e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.8915 $Y=0.1590 $X2=0.8780 $Y2=0.1590
r35 18 19 7.66224 $w=2.02e-08 $l=1.3e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9045 $Y=0.1590 $X2=0.8915 $Y2=0.1590
r36 17 18 9.13575 $w=2.02e-08 $l=1.55e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9200 $Y=0.1590 $X2=0.9045 $Y2=0.1590
r37 16 17 9.13575 $w=2.02e-08 $l=1.55e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9355 $Y=0.1590 $X2=0.9200 $Y2=0.1590
r38 5 16 22.3973 $w=2.02e-08 $l=3.8e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9735 $Y=0.1590 $X2=0.9355 $Y2=0.1590
r39 3 15 3.13392 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.9990
+ $Y=0.1590 $X2=0.9990 $Y2=0.1590
r40 3 5 24.6471 $w=2.06454e-08 $l=2.55e-08 $layer=LISD $thickness=3.21959e-08
+ $X=0.9990 $Y=0.1590 $X2=0.9735 $Y2=0.1590
r41 9 15 0.314665 $w=2.27e-07 $l=2.4e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.9990 $Y=0.1350 $X2=0.9990 $Y2=0.1590
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%MS VSS 14 70 71 74 76 87 89 4 1 23 19 28 20
+ 22 16 25 5 24 21 3 27 15 18 17
c1 1 VSS 0.000889461f
c2 3 VSS 0.00795946f
c3 4 VSS 0.00878592f
c4 5 VSS 0.00928199f
c5 14 VSS 0.032781f
c6 15 VSS 0.00351867f
c7 16 VSS 0.00229424f
c8 17 VSS 0.00277688f
c9 18 VSS 0.00270789f
c10 19 VSS 0.0022832f
c11 20 VSS 0.000655584f
c12 21 VSS 0.00961029f
c13 22 VSS 0.00238124f
c14 23 VSS 0.00480972f
c15 24 VSS 0.00321907f
c16 25 VSS 0.00220474f
c17 26 VSS 0.00134658f
c18 27 VSS 0.00601192f
c19 28 VSS 0.0077478f
r1 16 84 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9035 $Y=0.0405 $X2=0.9160 $Y2=0.0405
r2 89 16 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9010 $Y=0.0405 $X2=0.9035 $Y2=0.0405
r3 87 86 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9890 $Y=0.0405 $X2=0.9865 $Y2=0.0405
r4 17 86 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9740 $Y=0.0405 $X2=0.9865 $Y2=0.0405
r5 84 85 6.58477 $w=2.32e-08 $l=1.4e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.9180 $Y=0.0405 $X2=0.9320 $Y2=0.0405
r6 5 17 11.7585 $w=2.32e-08 $l=2.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.9470
+ $Y=0.0405 $X2=0.9720 $Y2=0.0405
r7 5 85 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.9470
+ $Y=0.0405 $X2=0.9320 $Y2=0.0405
r8 82 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.9720 $Y=0.0450
+ $X2=0.9720 $Y2=0.0405
r9 81 82 7.81186 $w=1.3e-08 $l=3.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.9720
+ $Y=0.0785 $X2=0.9720 $Y2=0.0450
r10 80 81 13.2918 $w=1.3e-08 $l=5.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.9720
+ $Y=0.1355 $X2=0.9720 $Y2=0.0785
r11 24 27 6.51495 $w=1.43636e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9720 $Y=0.1920 $X2=0.9720 $Y2=0.2250
r12 24 80 13.1752 $w=1.3e-08 $l=5.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.9720
+ $Y=0.1920 $X2=0.9720 $Y2=0.1355
r13 77 78 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.9830
+ $Y=0.2250 $X2=0.9940 $Y2=0.2250
r14 27 77 1.38478 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9720 $Y=0.2250 $X2=0.9830 $Y2=0.2250
r15 76 75 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8270 $Y=0.2295 $X2=0.8245 $Y2=0.2295
r16 19 75 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8120 $Y=0.2295 $X2=0.8245 $Y2=0.2295
r17 72 73 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7415 $Y=0.2160 $X2=0.7460 $Y2=0.2160
r18 74 72 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.2160 $X2=0.7415 $Y2=0.2160
r19 18 73 0.185185 $w=5.4e-08 $l=1e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7560 $Y=0.2160 $X2=0.7460 $Y2=0.2160
r20 71 69 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.0405 $X2=0.7165 $Y2=0.0405
r21 3 69 0.537037 $w=2.7e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7020 $Y=0.0405 $X2=0.7165 $Y2=0.0405
r22 15 3 0.537037 $w=2.7e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.0405 $X2=0.7020 $Y2=0.0405
r23 70 15 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.0405 $X2=0.6875 $Y2=0.0405
r24 66 78 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.9940 $Y=0.2250
+ $X2=0.9940 $Y2=0.2250
r25 65 66 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M2 $thickness=3.6e-08 $X=0.9555
+ $Y=0.2250 $X2=0.9940 $Y2=0.2250
r26 64 65 25.7675 $w=1.3e-08 $l=1.105e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.8450 $Y=0.2250 $X2=0.9555 $Y2=0.2250
r27 63 64 20.9871 $w=1.3e-08 $l=9e-08 $layer=M2 $thickness=3.6e-08 $X=0.7550
+ $Y=0.2250 $X2=0.8450 $Y2=0.2250
r28 28 63 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.7435
+ $Y=0.2250 $X2=0.7550 $Y2=0.2250
r29 61 19 4.04632 $w=5.02e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7830 $Y=0.2160 $X2=0.8100 $Y2=0.2160
r30 4 61 4.04632 $w=5.02e-08 $l=2.7e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7560 $Y=0.2160 $X2=0.7830 $Y2=0.2160
r31 4 57 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7560 $Y=0.2160
+ $X2=0.7560 $Y2=0.2250
r32 59 60 7.95695 $w=2.02e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7020 $Y=0.0585 $X2=0.7020 $Y2=0.0720
r33 3 59 10.6093 $w=2.02e-08 $l=1.8e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7020 $Y=0.0405 $X2=0.7020 $Y2=0.0585
r34 57 63 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.7560 $Y=0.2250
+ $X2=0.7550 $Y2=0.2250
r35 56 57 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.7465
+ $Y=0.2250 $X2=0.7560 $Y2=0.2250
r36 55 56 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.7375
+ $Y=0.2250 $X2=0.7465 $Y2=0.2250
r37 23 26 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7200
+ $Y=0.2250 $X2=0.7020 $Y2=0.2250
r38 23 55 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.7200
+ $Y=0.2250 $X2=0.7375 $Y2=0.2250
r39 50 51 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.0765 $X2=0.7020 $Y2=0.0855
r40 50 60 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7020 $Y=0.0765
+ $X2=0.7020 $Y2=0.0720
r41 49 51 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.0990 $X2=0.7020 $Y2=0.0855
r42 48 49 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.1170 $X2=0.7020 $Y2=0.0990
r43 47 48 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.1295 $X2=0.7020 $Y2=0.1170
r44 46 47 5.47996 $w=1.3e-08 $l=2.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.1530 $X2=0.7020 $Y2=0.1295
r45 45 46 5.47996 $w=1.3e-08 $l=2.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.1765 $X2=0.7020 $Y2=0.1530
r46 44 45 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.1890 $X2=0.7020 $Y2=0.1765
r47 43 44 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.2005 $X2=0.7020 $Y2=0.1890
r48 22 26 2.43413 $w=1.59032e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7020 $Y=0.2095 $X2=0.7020 $Y2=0.2250
r49 22 43 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.2095 $X2=0.7020 $Y2=0.2005
r50 26 42 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7020 $Y=0.2250 $X2=0.6805 $Y2=0.2250
r51 41 42 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.6400
+ $Y=0.2250 $X2=0.6805 $Y2=0.2250
r52 40 41 6.99569 $w=1.3e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.6100
+ $Y=0.2250 $X2=0.6400 $Y2=0.2250
r53 21 25 4.19024 $w=1.40976e-08 $l=2.54018e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5920 $Y=0.2250 $X2=0.5670 $Y2=0.2205
r54 21 40 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5920
+ $Y=0.2250 $X2=0.6100 $Y2=0.2250
r55 25 38 2.55791 $w=1.46667e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.2205 $X2=0.5670 $Y2=0.2070
r56 37 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1935 $X2=0.5670 $Y2=0.2070
r57 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1800 $X2=0.5670 $Y2=0.1935
r58 20 36 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1675 $X2=0.5670 $Y2=0.1800
r59 1 32 5.31651 $w=1.53e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.5670
+ $Y=0.1800 $X2=0.5670 $Y2=0.1800
r60 1 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1800
+ $X2=0.5670 $Y2=0.1800
r61 14 32 0.314665 $w=2.27e-07 $l=4.5e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5670 $Y=0.1350 $X2=0.5670 $Y2=0.1800
r62 4 18 1e-05
.ends

.subckt PM_ASYNC_DFFHx1_ASAP7_75t_R%CLKB VSS 11 12 69 71 20 15 5 6 18 19 17 13
+ 14 1 16 2
c1 1 VSS 0.000142521f
c2 2 VSS 9.70139e-20
c3 5 VSS 0.00737785f
c4 6 VSS 0.00695769f
c5 11 VSS 0.00448265f
c6 12 VSS 0.00493822f
c7 13 VSS 0.00643627f
c8 14 VSS 0.0063635f
c9 15 VSS 0.00335405f
c10 16 VSS 0.000965112f
c11 17 VSS 0.00128187f
c12 18 VSS 0.00631154f
c13 19 VSS 0.00547758f
c14 20 VSS 0.021422f
r1 14 6 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1600 $Y2=0.2160
r2 71 14 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r3 13 5 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1600 $Y2=0.0540
r4 69 13 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r5 6 61 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1655 $Y2=0.2340
r6 5 57 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1655 $Y2=0.0360
r7 1 55 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
r8 11 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r9 61 62 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1655
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r10 19 51 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2340 $X2=0.1890 $Y2=0.2125
r11 19 62 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2340 $X2=0.1755 $Y2=0.2340
r12 57 58 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1655
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r13 18 48 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1890 $Y2=0.0575
r14 18 58 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1755 $Y2=0.0360
r15 55 56 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1555
r16 16 52 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1735 $X2=0.4050 $Y2=0.1890
r17 16 56 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1735 $X2=0.4050 $Y2=0.1555
r18 50 51 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1990 $X2=0.1890 $Y2=0.2125
r19 49 50 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1900 $X2=0.1890 $Y2=0.1990
r20 47 48 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0790 $X2=0.1890 $Y2=0.0575
r21 46 47 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0970 $X2=0.1890 $Y2=0.0790
r22 45 46 9.211 $w=1.3e-08 $l=3.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1365 $X2=0.1890 $Y2=0.0970
r23 44 49 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1810 $X2=0.1890 $Y2=0.1900
r24 15 44 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1735 $X2=0.1890 $Y2=0.1810
r25 15 45 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1735 $X2=0.1890 $Y2=0.1365
r26 41 42 40.2252 $w=1.3e-08 $l=1.725e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.4050 $Y=0.1890 $X2=0.5775 $Y2=0.1890
r27 41 52 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4050 $Y=0.1890
+ $X2=0.4050 $Y2=0.1890
r28 40 41 25.1845 $w=1.3e-08 $l=1.08e-07 $layer=M2 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1890 $X2=0.4050 $Y2=0.1890
r29 39 40 25.1845 $w=1.3e-08 $l=1.08e-07 $layer=M2 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1890 $X2=0.2970 $Y2=0.1890
r30 39 49 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1890 $Y=0.1890
+ $X2=0.1890 $Y2=0.1900
r31 37 42 51.0686 $w=1.3e-08 $l=2.19e-07 $layer=M2 $thickness=3.6e-08 $X=0.7965
+ $Y=0.1890 $X2=0.5775 $Y2=0.1890
r32 20 35 5.59655 $w=1.3e-08 $l=2.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.8670
+ $Y=0.1890 $X2=0.8910 $Y2=0.1890
r33 20 37 16.4399 $w=1.3e-08 $l=7.05e-08 $layer=M2 $thickness=3.6e-08 $X=0.8670
+ $Y=0.1890 $X2=0.7965 $Y2=0.1890
r34 33 35 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.8910 $Y=0.1890
+ $X2=0.8910 $Y2=0.1890
r35 32 33 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1765 $X2=0.8910 $Y2=0.1890
r36 31 32 1.51573 $w=1.3e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1700 $X2=0.8910 $Y2=0.1765
r37 30 31 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1435 $X2=0.8910 $Y2=0.1700
r38 29 30 7.57867 $w=1.3e-08 $l=3.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1110 $X2=0.8910 $Y2=0.1435
r39 28 29 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1005 $X2=0.8910 $Y2=0.1110
r40 17 28 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.0980 $X2=0.8910 $Y2=0.1005
r41 2 25 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.8910
+ $Y=0.1110 $X2=0.8910 $Y2=0.1110
r42 2 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8910 $Y=0.1110
+ $X2=0.8910 $Y2=0.1110
r43 12 25 0.314665 $w=2.27e-07 $l=2.4e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.8910 $Y=0.1350 $X2=0.8910 $Y2=0.1110
.ends


*
.SUBCKT ASYNC_DFFHx1_ASAP7_75t_R VSS VDD CLK D RESET SET QN
*
* VSS VSS
* VDD VDD
* CLK CLK
* D D
* RESET RESET
* SET SET
* QN QN
*
*

MM20 N_MM20_d N_MM20_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM23 N_MM23_d N_MM22_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM1_g N_MM9_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM48 N_MM48_d N_MM49_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM47 N_MM47_d N_MM46_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM6 N_MM6_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM43 N_MM43_d N_MM43_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM34 N_MM34_d N_MM34_g N_MM34_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM12 N_MM12_d N_MM12_g N_MM12_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM47@2 N_MM47@2_d N_MM47@2_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM44 N_MM44_d N_MM44_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM29 N_MM29_d N_MM29_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM33 N_MM33_d N_MM33_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM24 N_MM24_d N_MM24_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM21 N_MM21_d N_MM20_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM22 N_MM22_d N_MM22_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM11 N_MM11_d N_MM11_g N_MM11_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM49 N_MM49_d N_MM49_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM46 N_MM46_d N_MM46_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM7 N_MM7_d N_MM7_g N_MM7_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM13 N_MM13_d N_MM34_g N_MM13_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM35 N_MM35_d N_MM12_g N_MM35_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM37 N_MM37_d N_MM37_g N_MM37_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM42 N_MM42_d N_MM47@2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM45 N_MM45_d N_MM44_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM28 N_MM28_d N_MM29_g N_MM28_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM25 N_MM25_d N_MM24_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "ASYNC_DFFHx1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "ASYNC_DFFHx1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%NET077 VSS N_MM37_s N_MM42_d N_NET077_1
+ PM_ASYNC_DFFHx1_ASAP7_75t_R%NET077
cc_1 N_NET077_1 N_MM47@2_g 0.0127072f
cc_2 N_NET077_1 N_MM37_g 0.012521f
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_ASYNC_DFFHx1_ASAP7_75t_R%noxref_24
cc_3 N_noxref_24_1 N_MM20_g 0.00832651f
cc_4 N_noxref_24_1 N_CLKN_30 6.65464e-20
cc_5 N_noxref_24_1 N_CLKN_29 6.97178e-20
cc_6 N_noxref_24_1 N_CLKN_27 7.17979e-20
cc_7 N_noxref_24_1 N_CLKN_28 0.00013996f
cc_8 N_noxref_24_1 N_CLKN_22 0.000255836f
cc_9 N_noxref_24_1 N_CLKN_21 0.000465584f
cc_10 N_noxref_24_1 N_CLKN_10 0.000485078f
cc_11 N_noxref_24_1 N_CLKN_9 0.000566938f
cc_12 N_noxref_24_1 N_CLKN_19 0.0129306f
cc_13 N_noxref_24_1 N_CLKN_20 0.0423165f
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%PD1 VSS N_MM5_d N_MM4_s N_PD1_1
+ PM_ASYNC_DFFHx1_ASAP7_75t_R%PD1
cc_14 N_PD1_1 N_MM4_g 0.0170489f
cc_15 N_PD1_1 N_MM3_g 0.0170754f
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_ASYNC_DFFHx1_ASAP7_75t_R%noxref_25
cc_16 N_noxref_25_1 N_MM22_g 0.0033982f
cc_17 N_noxref_25_1 N_CLKN_1 0.00557704f
cc_18 N_noxref_25_1 N_CLKB_15 0.000297581f
cc_19 N_noxref_25_1 N_CLKB_6 0.000449073f
cc_20 N_noxref_25_1 N_CLKB_5 0.000450808f
cc_21 N_noxref_25_1 N_CLKB_13 0.0128254f
cc_22 N_noxref_25_1 N_CLKB_14 0.0412445f
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%CLK VSS CLK N_MM20_g N_CLK_8 N_CLK_5 N_CLK_1
+ N_CLK_6 N_CLK_4 N_CLK_7 PM_ASYNC_DFFHx1_ASAP7_75t_R%CLK
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%noxref_26 VSS N_noxref_26_1
+ PM_ASYNC_DFFHx1_ASAP7_75t_R%noxref_26
cc_23 N_noxref_26_1 N_D_1 0.00462337f
cc_24 N_noxref_26_1 N_CLKB_5 0.000111851f
cc_25 N_noxref_26_1 N_CLKB_15 0.000194781f
cc_26 N_noxref_26_1 N_CLKB_14 0.000993265f
cc_27 N_noxref_26_1 N_noxref_25_1 0.0181393f
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%D VSS D N_MM3_g N_D_6 N_D_4 N_D_1 N_D_5 N_D_8
+ N_D_9 PM_ASYNC_DFFHx1_ASAP7_75t_R%D
cc_28 N_MM3_g N_CLKN_23 8.04196e-20
cc_29 N_MM3_g N_CLKN_1 0.000100561f
cc_30 N_MM3_g N_CLKN_30 0.000410223f
cc_31 N_MM3_g N_CLKN_24 0.00025369f
cc_32 N_MM3_g N_CLKN_2 0.000593503f
cc_33 N_D_6 N_CLKN_24 0.000574098f
cc_34 N_D_4 N_CLKN_30 0.000630478f
cc_35 N_D_6 N_CLKN_30 0.000926088f
cc_36 N_D_1 N_CLKN_2 0.00134023f
cc_37 N_D_5 N_CLKN_30 0.00231994f
cc_38 N_MM3_g N_MM4_g 0.0053599f
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%NET078 VSS N_MM11_s N_MM49_d N_NET078_1
+ PM_ASYNC_DFFHx1_ASAP7_75t_R%NET078
cc_39 N_NET078_1 N_MM11_g 0.00779128f
cc_40 N_NET078_1 N_MM49_g 0.00779979f
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%PD2 VSS N_MM35_s N_MM37_d N_PD2_1
+ PM_ASYNC_DFFHx1_ASAP7_75t_R%PD2
cc_41 N_PD2_1 N_MM12_g 0.0125496f
cc_42 N_PD2_1 N_SH_16 0.000305942f
cc_43 N_PD2_1 N_MM37_g 0.0126785f
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%NET076 VSS N_MM45_d N_MM28_s N_NET076_1
+ PM_ASYNC_DFFHx1_ASAP7_75t_R%NET076
cc_44 N_NET076_1 N_MM44_g 0.0125534f
cc_45 N_NET076_1 N_MM29_g 0.0125943f
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%noxref_29 VSS N_noxref_29_1
+ PM_ASYNC_DFFHx1_ASAP7_75t_R%noxref_29
cc_46 N_noxref_29_1 N_MM24_g 0.00398669f
cc_47 N_noxref_29_1 N_noxref_28_1 0.018422f
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%noxref_30 VSS N_noxref_30_1
+ PM_ASYNC_DFFHx1_ASAP7_75t_R%noxref_30
cc_48 N_noxref_30_1 N_MM24_g 0.00379402f
cc_49 N_noxref_30_1 N_QN_7 0.0172859f
cc_50 N_noxref_30_1 N_QN_8 0.0611488f
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%QN VSS QN N_MM24_d N_MM25_d N_QN_7 N_QN_2 N_QN_1
+ N_QN_8 N_QN_9 PM_ASYNC_DFFHx1_ASAP7_75t_R%QN
cc_51 N_QN_7 N_SH_21 0.00127234f
cc_52 N_QN_7 N_SH_2 0.000796123f
cc_53 N_QN_7 N_SH_23 0.000958532f
cc_54 N_QN_2 N_MM24_g 0.00119368f
cc_55 N_QN_1 N_MM24_g 0.00126944f
cc_56 N_QN_8 N_SH_2 0.00185919f
cc_57 N_QN_8 N_MM24_g 0.0151479f
cc_58 N_QN_9 N_SH_21 0.00551344f
cc_59 N_QN_7 N_MM24_g 0.0544374f
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%SS VSS N_MM37_g N_MM33_g N_MM28_d N_MM44_d
+ N_MM29_d N_SS_3 N_SS_15 N_SS_4 N_SS_7 N_SS_9 N_SS_1 N_SS_16 N_SS_6 N_SS_8
+ N_SS_5 PM_ASYNC_DFFHx1_ASAP7_75t_R%SS
cc_60 N_MM37_g N_CLKB_2 0.000529903f
cc_61 N_SS_3 N_CLKB_2 0.00121116f
cc_62 N_MM37_g N_MM12_g 0.0102985f
cc_63 N_MM37_g N_MS_5 0.00222406f
cc_64 N_MM37_g N_MS_16 0.00752934f
cc_65 N_SS_3 N_MS_24 0.00126022f
cc_66 N_SS_3 N_MS_17 0.00261353f
cc_67 N_MM37_g N_MS_17 0.0242126f
cc_68 N_SS_15 N_MM44_g 0.00674774f
cc_69 N_SS_4 N_MM44_g 0.000524025f
cc_70 N_SS_3 N_RESET_2 0.0025198f
cc_71 N_SS_3 N_RESET_9 0.000720208f
cc_72 N_SS_7 N_RESET_2 0.00100414f
cc_73 N_SS_3 N_MM44_g 0.0141085f
cc_74 N_SS_3 N_MM47@2_g 0.00306439f
cc_75 N_MM37_g N_SET_5 0.0030766f
cc_76 N_MM37_g N_MM47@2_g 0.0144679f
cc_77 N_MM33_g N_SH_21 7.65444e-20
cc_78 N_MM33_g N_SH_20 8.45622e-20
cc_79 N_SS_15 N_MM29_g 0.00677165f
cc_80 N_SS_9 N_SH_1 0.00028751f
cc_81 N_SS_1 N_SH_19 0.000314665f
cc_82 N_SS_16 N_MM29_g 0.0112505f
cc_83 N_SS_6 N_SH_23 0.000521059f
cc_84 N_SS_4 N_MM29_g 0.000531037f
cc_85 N_SS_8 N_MM29_g 0.000912145f
cc_86 N_SS_5 N_SH_1 0.00617288f
cc_87 N_SS_7 N_SH_1 0.000995867f
cc_88 N_SS_5 N_SH_20 0.00126239f
cc_89 N_SS_3 N_SH_19 0.00134184f
cc_90 N_SS_6 N_SH_1 0.00190844f
cc_91 N_MM37_g N_SH_6 0.00203159f
cc_92 N_MM33_g N_MM29_g 0.0334749f
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%noxref_28 VSS N_noxref_28_1
+ PM_ASYNC_DFFHx1_ASAP7_75t_R%noxref_28
cc_93 N_noxref_28_1 N_MM24_g 0.00076718f
cc_94 N_noxref_28_1 N_SS_6 0.000782314f
cc_95 N_noxref_28_1 N_MM33_g 0.0167259f
cc_96 N_noxref_28_1 N_PD3_8 0.0166207f
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%SH VSS N_MM29_g N_MM24_g N_MM35_d N_MM13_s
+ N_MM34_d N_MM12_s N_SH_14 N_SH_5 N_SH_23 N_SH_15 N_SH_18 N_SH_17 N_SH_16
+ N_SH_7 N_SH_6 N_SH_19 N_SH_22 N_SH_1 N_SH_20 N_SH_21 N_SH_2
+ PM_ASYNC_DFFHx1_ASAP7_75t_R%SH
cc_97 N_SH_14 N_CLKN_30 0.000106253f
cc_98 N_SH_5 N_MM34_g 0.00088022f
cc_99 N_SH_23 N_CLKN_30 0.000126804f
cc_100 N_SH_15 N_MM34_g 0.00014475f
cc_101 N_SH_18 N_CLKN_26 0.000151251f
cc_102 N_SH_17 N_MM34_g 0.00016522f
cc_103 N_SH_5 N_CLKN_4 0.000264595f
cc_104 N_SH_16 N_MM34_g 0.0113919f
cc_105 N_SH_7 N_MM34_g 0.000301957f
cc_106 N_SH_5 N_CLKN_26 0.000433337f
cc_107 N_SH_14 N_CLKN_4 0.000646729f
cc_108 N_SH_14 N_MM34_g 0.0379585f
cc_109 N_SH_15 N_MM12_g 0.000167352f
cc_110 N_SH_14 N_MM12_g 0.0116478f
cc_111 N_SH_18 N_CLKB_17 0.0003012f
cc_112 N_SH_6 N_CLKB_17 0.000344996f
cc_113 N_SH_7 N_MM12_g 0.0003929f
cc_114 N_SH_19 N_CLKB_17 0.0110656f
cc_115 N_SH_14 N_CLKB_2 0.000798887f
cc_116 N_SH_5 N_MM12_g 0.000826391f
cc_117 N_SH_19 N_CLKB_2 0.000871405f
cc_118 N_SH_6 N_MM12_g 0.00132042f
cc_119 N_SH_23 N_CLKB_20 0.00154747f
cc_120 N_SH_7 N_CLKB_20 0.00168235f
cc_121 N_SH_16 N_MM12_g 0.0389532f
cc_122 N_SH_5 N_MS_24 0.000174163f
cc_123 N_SH_6 N_MS_24 0.00052448f
cc_124 N_SH_16 N_MS_19 0.000594762f
cc_125 N_SH_19 N_MS_27 0.000922882f
cc_126 N_SH_14 N_MS_16 0.000592156f
cc_127 N_SH_18 N_MS_5 0.00028709f
cc_128 N_SH_22 N_MS_5 0.00168728f
cc_129 N_SH_5 N_MS_5 0.000510395f
cc_130 N_SH_22 N_MS_24 0.000608397f
cc_131 N_SH_7 N_MS_4 0.000929482f
cc_132 N_SH_16 N_MS_4 0.000964689f
cc_133 N_SH_19 N_MS_28 0.00174538f
cc_134 N_SH_23 N_MS_28 0.00235516f
cc_135 N_SH_19 N_MS_24 0.00962132f
cc_136 N_SH_19 N_RESET_12 0.000741463f
cc_137 N_SH_23 N_RESET_9 0.000548544f
cc_138 N_SH_1 N_RESET_2 0.00246392f
cc_139 N_SH_20 N_RESET_9 0.00332037f
cc_140 N_MM29_g N_MM44_g 0.0104239f
cc_141 N_SH_23 N_RESET_12 0.0146435f
cc_142 N_SH_5 N_SET_5 8.32109e-20
cc_143 N_SH_14 N_SET_5 8.58551e-20
cc_144 N_SH_20 N_SET_12 0.000110751f
cc_145 N_SH_18 N_SET_11 0.000119938f
cc_146 N_MM29_g N_MM47@2_g 0.000202222f
cc_147 N_SH_18 N_SET_12 0.000319793f
cc_148 N_SH_6 N_SET_5 0.00298746f
cc_149 N_SH_23 N_SET_12 0.000464978f
cc_150 N_SH_7 N_SET_5 0.00100621f
cc_151 N_SH_19 N_SET_5 0.00123521f
cc_152 N_SH_19 N_SET_12 0.00128516f
cc_153 N_SH_16 N_SET_5 0.00548907f
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%NET079 VSS N_MM46_d N_MM7_s N_NET079_1
+ PM_ASYNC_DFFHx1_ASAP7_75t_R%NET079
cc_154 N_NET079_1 N_MM7_g 0.0126468f
cc_155 N_NET079_1 N_MM46_g 0.0125887f
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%NET051 VSS N_MM10_s N_MM11_d N_NET051_4
+ N_NET051_5 N_NET051_1 PM_ASYNC_DFFHx1_ASAP7_75t_R%NET051
cc_156 N_NET051_4 N_MM10_g 0.0152527f
cc_157 N_NET051_5 N_MS_20 0.000212383f
cc_158 N_NET051_1 N_MS_1 0.0003086f
cc_159 N_NET051_5 N_MS_1 0.000555691f
cc_160 N_NET051_1 N_MM11_g 0.0012459f
cc_161 N_NET051_5 N_MM11_g 0.0153141f
cc_162 N_NET051_1 N_MH_13 0.000301799f
cc_163 N_NET051_4 N_MH_13 0.000346228f
cc_164 N_NET051_1 N_MH_17 0.000585782f
cc_165 N_NET051_4 N_MH_4 0.000630192f
cc_166 N_NET051_1 N_MH_21 0.00238192f
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%RESET VSS RESET N_MM49_g N_MM44_g N_RESET_12
+ N_RESET_10 N_RESET_7 N_RESET_8 N_RESET_2 N_RESET_9 N_RESET_11 N_RESET_1
+ PM_ASYNC_DFFHx1_ASAP7_75t_R%RESET
cc_167 N_RESET_12 N_CLKN_26 0.000750984f
cc_168 N_RESET_10 N_CLKN_30 0.000297484f
cc_169 N_RESET_7 N_CLKN_30 0.000533286f
cc_170 N_RESET_12 N_CLKN_30 0.0179573f
cc_171 N_RESET_12 N_CLKB_20 0.00214826f
cc_172 N_RESET_8 N_CLKB_20 0.000387276f
cc_173 N_RESET_12 N_CLKB_17 0.00200404f
cc_174 N_MM49_g N_MS_24 9.43794e-20
cc_175 N_MM49_g N_MS_3 0.000203605f
cc_176 N_RESET_2 N_MS_24 0.000143922f
cc_177 N_RESET_9 N_MS_27 0.000169417f
cc_178 N_RESET_10 N_MS_22 0.00369577f
cc_179 N_RESET_10 N_MS_20 0.000231711f
cc_180 N_RESET_9 N_MS_24 0.000760037f
cc_181 N_RESET_7 N_MS_20 0.000799295f
cc_182 N_RESET_11 N_MS_20 0.000927275f
cc_183 N_RESET_1 N_MS_1 0.00271279f
cc_184 N_RESET_12 N_MS_24 0.00137344f
cc_185 N_RESET_11 N_MS_21 0.0014664f
cc_186 N_RESET_12 N_MS_28 0.00172657f
cc_187 N_RESET_8 N_MS_21 0.00511545f
cc_188 N_MM49_g N_MM11_g 0.0110456f
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%PU1 VSS N_MM3_d N_MM1_s N_PU1_5 N_PU1_4 N_PU1_1
+ PM_ASYNC_DFFHx1_ASAP7_75t_R%PU1
cc_189 N_PU1_5 N_CLKN_2 0.00205667f
cc_190 N_PU1_5 N_CLKN_24 0.000545742f
cc_191 N_PU1_5 N_MM4_g 0.0738133f
cc_192 N_PU1_4 N_MM3_g 0.0358725f
cc_193 N_PU1_5 N_CLKB_1 0.000836281f
cc_194 N_PU1_5 N_CLKB_16 0.000665519f
cc_195 N_PU1_5 N_MM1_g 0.0348684f
cc_196 N_PU1_1 N_MH_4 0.0013618f
cc_197 N_PU1_1 N_MH_13 0.00295732f
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%NET020 VSS N_MM9_s N_MM8_d N_MM48_d N_NET020_7
+ N_NET020_1 N_NET020_8 N_NET020_2 N_NET020_9 PM_ASYNC_DFFHx1_ASAP7_75t_R%NET020
cc_198 N_NET020_7 N_CLKN_30 0.00011596f
cc_199 N_NET020_7 N_CLKN_3 0.000480358f
cc_200 N_NET020_7 N_CLKN_25 0.000509302f
cc_201 N_NET020_1 N_MM10_g 0.000738688f
cc_202 N_NET020_7 N_MM10_g 0.026327f
cc_203 N_NET020_7 N_CLKB_16 0.000165325f
cc_204 N_NET020_7 N_CLKB_1 0.000187051f
cc_205 N_NET020_7 N_MM1_g 0.0247033f
cc_206 N_NET020_8 N_MM11_g 0.0250462f
cc_207 N_NET020_8 N_RESET_10 0.000427811f
cc_208 N_NET020_2 N_MM49_g 0.000594907f
cc_209 N_NET020_8 N_MM49_g 0.0249706f
cc_210 N_NET020_9 N_MH_3 0.000203208f
cc_211 N_NET020_9 N_MH_17 0.000290004f
cc_212 N_NET020_1 N_MH_3 0.00288006f
cc_213 N_NET020_7 N_MH_10 0.000461528f
cc_214 N_NET020_7 N_MH_11 0.000505866f
cc_215 N_NET020_9 N_MH_15 0.000572984f
cc_216 N_NET020_9 N_MH_20 0.000890654f
cc_217 N_NET020_9 N_MH_22 0.00165521f
cc_218 N_NET020_9 N_MH_18 0.00678266f
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%noxref_27 VSS N_noxref_27_1
+ PM_ASYNC_DFFHx1_ASAP7_75t_R%noxref_27
cc_219 N_noxref_27_1 N_CLKN_3 0.000401179f
cc_220 N_noxref_27_1 N_MM10_g 0.0152284f
cc_221 N_noxref_27_1 N_MM11_g 0.0101851f
cc_222 N_noxref_27_1 N_MH_17 0.000265606f
cc_223 N_noxref_27_1 N_MH_13 0.00085633f
cc_224 N_noxref_27_1 N_NET051_1 0.000743632f
cc_225 N_noxref_27_1 N_NET051_4 0.00705131f
cc_226 N_noxref_27_1 N_NET051_5 0.0240396f
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%CLKN VSS N_MM22_g N_MM4_g N_MM10_g N_MM34_g
+ N_MM20_d N_MM21_d N_CLKN_28 N_CLKN_10 N_CLKN_9 N_CLKN_20 N_CLKN_19 N_CLKN_1
+ N_CLKN_23 N_CLKN_22 N_CLKN_27 N_CLKN_29 N_CLKN_21 N_CLKN_30 N_CLKN_24
+ N_CLKN_2 N_CLKN_25 N_CLKN_26 N_CLKN_4 N_CLKN_3
+ PM_ASYNC_DFFHx1_ASAP7_75t_R%CLKN
cc_227 N_CLKN_28 N_MM20_g 0.000222492f
cc_228 N_CLKN_10 N_MM20_g 0.0011032f
cc_229 N_CLKN_9 N_MM20_g 0.00112998f
cc_230 N_CLKN_20 N_MM20_g 0.0110783f
cc_231 N_CLKN_19 N_MM20_g 0.0113756f
cc_232 N_CLKN_1 N_MM20_g 0.000397316f
cc_233 N_CLKN_23 N_MM20_g 0.000571637f
cc_234 N_CLKN_22 N_CLK_8 0.000803041f
cc_235 N_CLKN_27 N_CLK_5 0.000819345f
cc_236 N_CLKN_28 N_CLK_1 0.000862467f
cc_237 N_CLKN_29 N_CLK_6 0.000899886f
cc_238 N_CLKN_21 N_CLK_4 0.00151266f
cc_239 N_CLKN_30 N_CLK_8 0.00161009f
cc_240 N_CLKN_29 N_CLK_8 0.00199449f
cc_241 N_CLKN_27 N_CLK_7 0.00210914f
cc_242 N_CLKN_23 N_CLK_8 0.00211464f
cc_243 N_CLKN_1 N_CLK_1 0.0024079f
cc_244 N_CLKN_28 N_CLK_4 0.00468657f
cc_245 N_MM22_g N_MM20_g 0.0350707f
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%PD3 VSS N_MM43_d N_MM34_s N_MM33_d N_PD3_7
+ N_PD3_1 N_PD3_11 N_PD3_9 N_PD3_10 N_PD3_8 N_PD3_2
+ PM_ASYNC_DFFHx1_ASAP7_75t_R%PD3
cc_246 N_PD3_7 N_CLKN_26 0.000508414f
cc_247 N_PD3_7 N_CLKN_30 0.00011117f
cc_248 N_PD3_7 N_CLKN_4 0.000882637f
cc_249 N_PD3_1 N_MM34_g 0.000790549f
cc_250 N_PD3_7 N_MM34_g 0.0250438f
cc_251 N_PD3_11 N_MS_24 0.00173222f
cc_252 N_PD3_11 N_RESET_12 0.00210855f
cc_253 N_PD3_11 N_MH_1 0.000134249f
cc_254 N_PD3_11 N_MH_19 0.000143038f
cc_255 N_PD3_9 N_MH_19 0.000550291f
cc_256 N_PD3_11 N_MH_22 0.00146867f
cc_257 N_PD3_11 N_SET_11 0.000248326f
cc_258 N_PD3_11 N_MM43_g 0.000333695f
cc_259 N_PD3_1 N_MM43_g 0.000650159f
cc_260 N_PD3_9 N_SET_11 0.00465807f
cc_261 N_PD3_7 N_MM43_g 0.0245094f
cc_262 N_PD3_11 N_SET_12 0.0202791f
cc_263 N_PD3_11 N_SH_20 0.000782923f
cc_264 N_PD3_11 N_MM29_g 9.3022e-20
cc_265 N_PD3_11 N_SH_21 0.000136953f
cc_266 N_PD3_11 N_SH_19 0.000270205f
cc_267 N_PD3_9 N_SH_18 0.00028875f
cc_268 N_PD3_1 N_SH_5 0.00246063f
cc_269 N_PD3_10 N_SH_20 0.000371471f
cc_270 N_PD3_7 N_SH_14 0.000797008f
cc_271 N_PD3_11 N_SH_18 0.000964294f
cc_272 N_PD3_11 N_SH_23 0.00166364f
cc_273 N_PD3_11 N_SH_22 0.00339169f
cc_274 N_PD3_8 N_SS_9 0.000922874f
cc_275 N_PD3_8 N_SS_6 0.000275669f
cc_276 N_PD3_10 N_SS_9 0.000283172f
cc_277 N_PD3_11 N_SS_3 0.000299346f
cc_278 N_PD3_2 N_MM33_g 0.000503549f
cc_279 N_PD3_8 N_MM33_g 0.0154457f
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%MH VSS N_MM7_g N_MM4_d N_MM9_d N_MM1_d N_MM10_d
+ N_MH_13 N_MH_18 N_MH_1 N_MH_11 N_MH_15 N_MH_14 N_MH_10 N_MH_19 N_MH_16
+ N_MH_20 N_MH_3 N_MH_17 N_MH_4 N_MH_22 N_MH_21 PM_ASYNC_DFFHx1_ASAP7_75t_R%MH
cc_280 N_MH_13 N_MM34_g 5.37954e-20
cc_281 N_MH_13 N_MM4_g 5.95147e-20
cc_282 N_MH_18 N_CLKN_30 0.000139218f
cc_283 N_MH_1 N_CLKN_4 0.000157598f
cc_284 N_MH_11 N_MM4_g 0.0244746f
cc_285 N_MH_15 N_CLKN_24 0.00218169f
cc_286 N_MH_14 N_MM10_g 0.000175136f
cc_287 N_MH_10 N_MM4_g 0.0101305f
cc_288 N_MH_19 N_CLKN_30 0.000217286f
cc_289 N_MH_18 N_CLKN_25 0.000219798f
cc_290 N_MH_16 N_CLKN_25 0.000249754f
cc_291 N_MH_20 N_CLKN_25 0.000255623f
cc_292 N_MH_3 N_CLKN_24 0.000288955f
cc_293 N_MH_17 N_CLKN_25 0.00734964f
cc_294 N_MH_3 N_CLKN_2 0.000521243f
cc_295 N_MH_10 N_CLKN_2 0.000840038f
cc_296 N_MH_17 N_CLKN_3 0.000951849f
cc_297 N_MH_13 N_CLKN_3 0.00122088f
cc_298 N_MH_3 N_MM4_g 0.00123421f
cc_299 N_MH_4 N_MM10_g 0.0012415f
cc_300 N_MH_22 N_CLKN_30 0.00946846f
cc_301 N_MH_13 N_MM10_g 0.0363287f
cc_302 N_MH_13 N_CLKB_16 0.000117672f
cc_303 N_MH_14 N_MM1_g 0.000144496f
cc_304 N_MH_21 N_CLKB_20 0.000178942f
cc_305 N_MH_16 N_CLKB_16 0.00139448f
cc_306 N_MH_10 N_MM1_g 0.0104787f
cc_307 N_MH_4 N_CLKB_16 0.00231447f
cc_308 N_MH_3 N_CLKB_16 0.000221217f
cc_309 N_MH_11 N_MM1_g 0.00556137f
cc_310 N_MH_19 N_CLKB_20 0.000473324f
cc_311 N_MH_4 N_CLKB_1 0.000646737f
cc_312 N_MH_15 N_CLKB_16 0.000659369f
cc_313 N_MH_22 N_CLKB_20 0.000866832f
cc_314 N_MH_17 N_CLKB_20 0.000922441f
cc_315 N_MH_3 N_MM1_g 0.000963245f
cc_316 N_MH_4 N_MM1_g 0.00132361f
cc_317 N_MH_13 N_CLKB_1 0.00147031f
cc_318 N_MH_16 N_CLKB_20 0.0017011f
cc_319 N_MH_13 N_MM1_g 0.0530163f
cc_320 N_MH_21 N_MS_25 0.000168143f
cc_321 N_MH_18 N_MM11_g 0.000177306f
cc_322 N_MH_18 N_MS_20 0.00018301f
cc_323 N_MH_17 N_MS_1 0.000534082f
cc_324 N_MH_17 N_MS_25 0.00021372f
cc_325 N_MM7_g N_MS_15 0.00673709f
cc_326 N_MH_19 N_MS_22 0.00731804f
cc_327 N_MM7_g N_MS_4 0.000340022f
cc_328 N_MH_19 N_MS_3 0.000540641f
cc_329 N_MH_1 N_MS_22 0.000541126f
cc_330 N_MH_22 N_MS_20 0.000819017f
cc_331 N_MH_1 N_MS_3 0.00101197f
cc_332 N_MM7_g N_MS_3 0.00123422f
cc_333 N_MH_17 N_MS_20 0.00175916f
cc_334 N_MM7_g N_MS_18 0.0338153f
cc_335 N_MH_18 N_RESET_10 0.000220282f
cc_336 N_MH_19 N_RESET_12 0.000636323f
cc_337 N_MH_22 N_RESET_10 0.00101887f
cc_338 N_MH_22 N_RESET_12 0.0112382f
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%SET VSS SET N_MM46_g N_MM43_g N_MM47@2_g N_SET_12
+ N_SET_11 N_SET_5 N_SET_10 N_SET_1 N_SET_3 PM_ASYNC_DFFHx1_ASAP7_75t_R%SET
cc_339 N_MM43_g N_CLKN_26 0.000388067f
cc_340 N_SET_12 N_CLKN_26 0.000386958f
cc_341 N_SET_11 N_CLKN_26 0.000585929f
cc_342 N_SET_5 N_CLKN_30 0.000733023f
cc_343 N_SET_5 N_CLKN_4 0.00220211f
cc_344 N_SET_5 N_MM34_g 0.00362494f
cc_345 N_SET_10 N_CLKN_26 0.00406314f
cc_346 N_MM43_g N_MM34_g 0.0108097f
cc_347 N_SET_5 N_CLKB_17 0.00144155f
cc_348 N_SET_5 N_CLKB_2 0.00126397f
cc_349 N_SET_10 N_CLKB_20 0.000812513f
cc_350 N_SET_5 N_MM12_g 0.005467f
cc_351 N_MM43_g N_MS_24 9.06176e-20
cc_352 N_SET_1 N_MS_22 0.000103221f
cc_353 N_SET_5 N_MS_27 0.000136124f
cc_354 N_MM47@2_g N_MS_5 0.000143704f
cc_355 N_SET_5 N_MS_4 0.00690448f
cc_356 N_SET_10 N_MS_28 0.000204848f
cc_357 N_MM46_g N_MS_15 0.00674777f
cc_358 N_MM47@2_g N_MS_17 0.0148648f
cc_359 N_MM43_g N_MS_19 0.00739443f
cc_360 N_SET_10 N_MS_23 0.000402254f
cc_361 N_SET_12 N_MS_24 0.000758253f
cc_362 N_SET_10 N_MS_22 0.000797662f
cc_363 N_SET_5 N_MS_22 0.0015703f
cc_364 N_SET_5 N_MS_24 0.00180182f
cc_365 N_MM43_g N_MS_4 0.00462483f
cc_366 N_MM46_g N_MS_3 0.0094043f
cc_367 N_MM43_g N_MS_18 0.0354642f
cc_368 N_SET_5 N_RESET_12 0.00196631f
cc_369 N_SET_5 N_RESET_10 0.000228974f
cc_370 N_SET_11 N_RESET_12 0.000290247f
cc_371 N_SET_5 N_RESET_9 0.000335087f
cc_372 N_SET_12 N_RESET_9 0.000353943f
cc_373 N_SET_3 N_RESET_2 0.000401779f
cc_374 N_SET_10 N_RESET_12 0.000467642f
cc_375 N_SET_1 N_RESET_1 0.000510913f
cc_376 N_SET_5 N_RESET_2 0.000517691f
cc_377 N_SET_5 N_RESET_1 0.000606711f
cc_378 N_MM46_g N_MM49_g 0.00755887f
cc_379 N_MM47@2_g N_MM44_g 0.00920011f
cc_380 N_SET_12 N_RESET_12 0.0213676f
cc_381 N_SET_11 N_MH_19 0.000976429f
cc_382 N_SET_12 N_MH_22 0.000457098f
cc_383 N_SET_5 N_MH_22 0.000506112f
cc_384 N_SET_10 N_MH_1 0.00072201f
cc_385 N_SET_10 N_MH_19 0.00325199f
cc_386 N_MM46_g N_MM7_g 0.00513406f
cc_387 N_SET_5 N_MH_1 0.00613245f
cc_388 N_MM43_g N_MM7_g 0.0142658f
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%MS VSS N_MM11_g N_MM47_d N_MM6_d N_MM7_d N_MM13_d
+ N_MM47@2_d N_MM12_d N_MS_4 N_MS_1 N_MS_23 N_MS_19 N_MS_28 N_MS_20 N_MS_22
+ N_MS_16 N_MS_25 N_MS_5 N_MS_24 N_MS_21 N_MS_3 N_MS_27 N_MS_15 N_MS_18 N_MS_17
+ PM_ASYNC_DFFHx1_ASAP7_75t_R%MS
cc_389 N_MS_4 N_CLKN_3 0.000122524f
cc_390 N_MS_4 N_CLKN_26 0.000334146f
cc_391 N_MS_4 N_CLKN_30 5.65663e-20
cc_392 N_MS_1 N_CLKN_30 8.79855e-20
cc_393 N_MS_23 N_CLKN_30 9.5963e-20
cc_394 N_MS_1 N_MM10_g 0.000100661f
cc_395 N_MM11_g N_MM10_g 0.00020639f
cc_396 N_MS_19 N_MM34_g 0.0066067f
cc_397 N_MS_28 N_CLKN_30 0.000428677f
cc_398 N_MS_20 N_CLKN_30 0.000470812f
cc_399 N_MS_22 N_CLKN_30 0.00204276f
cc_400 N_MS_4 N_MM34_g 0.00922665f
cc_401 N_MS_4 N_MM12_g 0.000123364f
cc_402 N_MS_16 N_CLKB_2 0.000145911f
cc_403 N_MS_16 N_MM12_g 0.0149374f
cc_404 N_MS_25 N_CLKB_20 0.000264551f
cc_405 N_MS_23 N_CLKB_20 0.000729881f
cc_406 N_MS_28 N_CLKB_17 0.000311709f
cc_407 N_MS_5 N_MM12_g 0.000317504f
cc_408 N_MS_24 N_CLKB_17 0.000466257f
cc_409 N_MS_22 N_CLKB_20 0.000596289f
cc_410 N_MS_21 N_CLKB_20 0.000866327f
cc_411 N_MS_20 N_CLKB_20 0.00100193f
cc_412 N_MS_28 N_CLKB_20 0.018514f
x_PM_ASYNC_DFFHx1_ASAP7_75t_R%CLKB VSS N_MM1_g N_MM12_g N_MM23_d N_MM22_d
+ N_CLKB_20 N_CLKB_15 N_CLKB_5 N_CLKB_6 N_CLKB_18 N_CLKB_19 N_CLKB_17 N_CLKB_13
+ N_CLKB_14 N_CLKB_1 N_CLKB_16 N_CLKB_2 PM_ASYNC_DFFHx1_ASAP7_75t_R%CLKB
cc_413 N_CLKB_20 N_CLK_6 0.000124881f
cc_414 N_CLKB_15 N_CLK_6 0.000595591f
cc_415 N_CLKB_5 N_CLK_6 0.000348623f
cc_416 N_CLKB_6 N_CLK_6 0.000366091f
cc_417 N_CLKB_18 N_CLK_6 0.000368507f
cc_418 N_CLKB_18 N_CLK_5 0.00117646f
cc_419 N_CLKB_19 N_CLK_6 0.0020005f
cc_420 N_CLKB_20 N_MM22_g 0.000151304f
cc_421 N_CLKB_17 N_CLKN_30 0.000129359f
cc_422 N_CLKB_13 N_MM22_g 0.0386163f
cc_423 N_CLKB_14 N_MM22_g 0.0112881f
cc_424 N_CLKB_19 N_CLKN_23 0.000345969f
cc_425 N_CLKB_18 N_CLKN_23 0.000354534f
cc_426 N_CLKB_1 N_CLKN_2 0.000802518f
cc_427 N_CLKB_16 N_CLKN_30 0.000423068f
cc_428 N_CLKB_20 N_CLKN_25 0.000430515f
cc_429 N_CLKB_15 N_CLKN_23 0.00811758f
cc_430 N_CLKB_20 N_CLKN_26 0.000491638f
cc_431 N_CLKB_15 N_CLKN_30 0.0005953f
cc_432 N_CLKB_5 N_MM22_g 0.000655069f
cc_433 N_CLKB_20 N_CLKN_24 0.000667067f
cc_434 N_CLKB_6 N_MM22_g 0.000683495f
cc_435 N_CLKB_15 N_CLKN_1 0.000693119f
cc_436 N_CLKB_2 N_CLKN_4 0.00192126f
cc_437 N_CLKB_1 N_CLKN_3 0.00275f
cc_438 N_CLKB_16 N_CLKN_24 0.00119903f
cc_439 N_CLKB_14 N_CLKN_1 0.00123094f
cc_440 N_MM1_g N_MM4_g 0.00160961f
cc_441 N_CLKB_17 N_CLKN_26 0.00310323f
cc_442 N_CLKB_16 N_CLKN_25 0.00362212f
cc_443 N_MM1_g N_MM10_g 0.00699089f
cc_444 N_MM12_g N_MM34_g 0.00711952f
cc_445 N_CLKB_20 N_CLKN_30 0.054386f
cc_446 N_MM1_g N_D_8 0.000112693f
cc_447 N_CLKB_6 N_D_8 0.000114499f
cc_448 N_CLKB_5 N_D_8 0.000118096f
cc_449 N_CLKB_18 N_D_8 0.000803939f
cc_450 N_CLKB_19 N_D_9 0.00107656f
cc_451 N_CLKB_20 N_D_6 0.00145553f
cc_452 N_CLKB_15 N_D_4 0.0017222f
cc_453 N_CLKB_15 N_D_5 0.00238656f
cc_454 N_CLKB_15 N_D_8 0.00435554f
*END of ASYNC_DFFHx1_ASAP7_75t_R.pxi
.ENDS
** Design:	ICGx1_ASAP7_75t_R
* Created:	"Fri Aug 17 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "ICGx1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "ICGx1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_ICGx1_ASAP7_75t_R%NOS1 VSS 2 3 1
c1 1 VSS 0.000877566f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2160 $X2=0.1080 $Y2=0.2160
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2160 $X2=0.1080 $Y2=0.2160
.ends

.subckt PM_ICGx1_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.00478343f
.ends

.subckt PM_ICGx1_ASAP7_75t_R%SE VSS 8 3 1 4
c1 1 VSS 0.00624099f
c2 3 VSS 0.0829922f
c3 4 VSS 0.00446073f
r1 9 10 2.3902 $w=1.3e-08 $l=1.03e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1267 $X2=0.1350 $Y2=0.1370
r2 8 9 0.408082 $w=1.3e-08 $l=1.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1250 $X2=0.1350 $Y2=0.1267
r3 8 4 6.47102 $w=1.3e-08 $l=2.78e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1250 $X2=0.1350 $Y2=0.0972
r4 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r5 1 10 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1370
.ends

.subckt PM_ICGx1_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.0320309f
.ends

.subckt PM_ICGx1_ASAP7_75t_R%ENA VSS 8 3 1 4
c1 1 VSS 0.00210225f
c2 3 VSS 0.0329591f
c3 4 VSS 0.00993401f
r1 9 10 2.3902 $w=1.3e-08 $l=1.03e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1267 $X2=0.0810 $Y2=0.1370
r2 8 9 0.408082 $w=1.3e-08 $l=1.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1250 $X2=0.0810 $Y2=0.1267
r3 8 4 6.47102 $w=1.3e-08 $l=2.78e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1250 $X2=0.0810 $Y2=0.0972
r4 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r5 1 10 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1370
.ends

.subckt PM_ICGx1_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.00458186f
.ends

.subckt PM_ICGx1_ASAP7_75t_R%noxref_26 VSS 1
c1 1 VSS 0.00481573f
.ends

.subckt PM_ICGx1_ASAP7_75t_R%GCLK VSS 20 15 25 7 9 1 2 8 10 11
c1 1 VSS 0.00805143f
c2 2 VSS 0.00816293f
c3 7 VSS 0.00371137f
c4 8 VSS 0.00376937f
c5 9 VSS 0.00603617f
c6 10 VSS 0.00387986f
c7 11 VSS 0.00336574f
c8 12 VSS 0.00290217f
c9 13 VSS 0.00321771f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9035 $Y=0.2025 $X2=0.9160 $Y2=0.2025
r2 25 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9010 $Y=0.2025 $X2=0.9035 $Y2=0.2025
r3 2 10 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.9180 $Y=0.2025
+ $X2=0.9180 $Y2=0.2340
r4 10 13 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9180 $Y=0.2340 $X2=0.9450 $Y2=0.2340
r5 13 22 2.6649 $w=1.77676e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.2340 $X2=0.9450 $Y2=0.2155
r6 21 22 6.8208 $w=1.3e-08 $l=2.93e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1862 $X2=0.9450 $Y2=0.2155
r7 20 21 4.72209 $w=1.3e-08 $l=2.02e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1660 $X2=0.9450 $Y2=0.1862
r8 20 19 12.0676 $w=1.3e-08 $l=5.18e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.1660 $X2=0.9450 $Y2=0.1142
r9 11 12 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.0540 $X2=0.9450 $Y2=0.0360
r10 11 19 14.0497 $w=1.3e-08 $l=6.02e-08 $layer=M1 $thickness=3.6e-08 $X=0.9450
+ $Y=0.0540 $X2=0.9450 $Y2=0.1142
r11 12 17 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9450 $Y=0.0360 $X2=0.9315 $Y2=0.0360
r12 16 17 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.0360 $X2=0.9315 $Y2=0.0360
r13 9 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.9045
+ $Y=0.0360 $X2=0.9180 $Y2=0.0360
r14 1 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.9180 $Y=0.0675
+ $X2=0.9180 $Y2=0.0360
r15 7 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9035 $Y=0.0675 $X2=0.9160 $Y2=0.0675
r16 15 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9010 $Y=0.0675 $X2=0.9035 $Y2=0.0675
.ends

.subckt PM_ICGx1_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.00423453f
.ends

.subckt PM_ICGx1_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.00439869f
.ends

.subckt PM_ICGx1_ASAP7_75t_R%NET0121 VSS 9 40 41 43 11 13 4 3 12 10 1 14
c1 1 VSS 0.00377593f
c2 3 VSS 0.00720448f
c3 4 VSS 0.00903034f
c4 9 VSS 0.0801794f
c5 10 VSS 0.0064067f
c6 11 VSS 0.00507154f
c7 12 VSS 0.016911f
c8 13 VSS 0.0107904f
c9 14 VSS 0.00655582f
c10 15 VSS 0.00372186f
c11 16 VSS 0.00354213f
r1 43 42 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r2 11 42 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r3 41 39 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0540 $X2=0.1225 $Y2=0.0540
r4 4 39 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0540 $X2=0.1225 $Y2=0.0540
r5 10 4 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0540 $X2=0.1080 $Y2=0.0540
r6 40 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0540 $X2=0.0935 $Y2=0.0540
r7 3 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0540 $Y2=0.2330
r8 4 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0540
+ $X2=0.1080 $Y2=0.0360
r9 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2330 $X2=0.0675 $Y2=0.2330
r10 34 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.2330 $X2=0.0675 $Y2=0.2330
r11 33 34 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2330 $X2=0.0810 $Y2=0.2330
r12 32 33 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2330 $X2=0.1080 $Y2=0.2330
r13 12 16 5.06479 $w=1.46038e-08 $l=2.70046e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1620 $Y=0.2330 $X2=0.1890 $Y2=0.2325
r14 12 32 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2330 $X2=0.1350 $Y2=0.2330
r15 29 30 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.1215 $Y2=0.0360
r16 27 30 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1215 $Y2=0.0360
r17 13 15 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1620 $Y=0.0360 $X2=0.1890 $Y2=0.0360
r18 13 27 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r19 16 25 0.983973 $w=1.77222e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2325 $X2=0.1890 $Y2=0.2235
r20 15 20 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1890 $Y2=0.0575
r21 24 25 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2110 $X2=0.1890 $Y2=0.2235
r22 23 24 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1985 $X2=0.1890 $Y2=0.2110
r23 22 23 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1910 $X2=0.1890 $Y2=0.1985
r24 21 22 9.211 $w=1.3e-08 $l=3.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1515 $X2=0.1890 $Y2=0.1910
r25 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0710 $X2=0.1890 $Y2=0.0575
r26 14 19 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0955 $X2=0.1890 $Y2=0.0710
r27 14 21 13.0586 $w=1.3e-08 $l=5.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0955 $X2=0.1890 $Y2=0.1515
r28 9 1 6.2219 $w=1.2115e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1340
r29 1 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1340
+ $X2=0.1890 $Y2=0.1515
r30 3 11 1e-05
.ends

.subckt PM_ICGx1_ASAP7_75t_R%PD1 VSS 7 10 4 5 1
c1 1 VSS 0.00996545f
c2 4 VSS 0.00323613f
c3 5 VSS 0.00185849f
r1 10 9 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r2 8 9 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2800 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r3 5 8 0.123457 $w=8.1e-08 $l=1e-08 $layer=N_src_drn $thickness=1e-09 $X=0.2700
+ $Y=0.0675 $X2=0.2800 $Y2=0.0675
r4 4 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0675 $X2=0.2140 $Y2=0.0675
r5 7 4 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2015 $Y2=0.0675
r6 1 5 1e-05
.ends

.subckt PM_ICGx1_ASAP7_75t_R%NET0140 VSS 2 3 1
c1 1 VSS 0.000863546f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.0675 $X2=0.7020 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.0675 $X2=0.7020 $Y2=0.0675
.ends

.subckt PM_ICGx1_ASAP7_75t_R%PU1 VSS 5 8 3 1
c1 1 VSS 0.00536668f
c2 3 VSS 0.00340271f
r1 8 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r2 6 7 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2260 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r3 1 6 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2140 $Y=0.2025 $X2=0.2260 $Y2=0.2025
r4 3 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2140 $Y2=0.2025
r5 5 3 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
.ends

.subckt PM_ICGx1_ASAP7_75t_R%PD3 VSS 5 8 3 1
c1 1 VSS 0.00335597f
c2 3 VSS 0.0024702f
r1 8 7 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0405 $X2=0.3925 $Y2=0.0405
r2 1 7 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3800 $Y=0.0405 $X2=0.3925 $Y2=0.0405
r3 4 1 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3680 $Y=0.0405 $X2=0.3800 $Y2=0.0405
r4 3 4 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.0405 $X2=0.3680 $Y2=0.0405
r5 5 3 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0405 $X2=0.3635 $Y2=0.0405
.ends

.subckt PM_ICGx1_ASAP7_75t_R%NET0141 VSS 2 3 1
c1 1 VSS 0.000908898f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.0675 $X2=0.8100 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8270 $Y=0.0675 $X2=0.8100 $Y2=0.0675
.ends

.subckt PM_ICGx1_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.00366369f
.ends

.subckt PM_ICGx1_ASAP7_75t_R%MS VSS 9 40 46 1 12 13 15 3 14 4 11 10
c1 1 VSS 0.00207698f
c2 3 VSS 0.00503664f
c3 4 VSS 0.0060406f
c4 9 VSS 0.0369206f
c5 10 VSS 0.00306582f
c6 11 VSS 0.00310462f
c7 12 VSS 0.00122337f
c8 13 VSS 0.0012459f
c9 14 VSS 0.00665905f
c10 15 VSS 0.000349358f
r1 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2295 $X2=0.4840 $Y2=0.2295
r2 46 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2295 $X2=0.4715 $Y2=0.2295
r3 4 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2295
+ $X2=0.4860 $Y2=0.2330
r4 42 43 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.2330 $X2=0.4990 $Y2=0.2330
r5 14 38 1.06916 $w=1.78e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.2330 $X2=0.5125 $Y2=0.2235
r6 14 43 1.90218 $w=1.65185e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5125 $Y=0.2330 $X2=0.4990 $Y2=0.2330
r7 10 31 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0405 $X2=0.4840 $Y2=0.0405
r8 40 10 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0405 $X2=0.4715 $Y2=0.0405
r9 37 38 2.49333 $w=1.4e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.2110 $X2=0.5125 $Y2=0.2235
r10 36 37 4.1888 $w=1.4e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.1900 $X2=0.5125 $Y2=0.2110
r11 35 36 3.69013 $w=1.4e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.1715 $X2=0.5125 $Y2=0.1900
r12 34 35 3.69013 $w=1.4e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.1530 $X2=0.5125 $Y2=0.1715
r13 33 34 4.1888 $w=1.4e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.1320 $X2=0.5125 $Y2=0.1530
r14 32 33 4.88693 $w=1.4e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.1075 $X2=0.5125 $Y2=0.1320
r15 13 15 0.843012 $w=1.80909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5125 $Y=0.0930 $X2=0.5125 $Y2=0.0820
r16 13 32 2.89227 $w=1.4e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.0930 $X2=0.5125 $Y2=0.1075
r17 3 29 10.904 $w=2.02e-08 $l=1.85e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4860 $Y=0.0635 $X2=0.4860 $Y2=0.0820
r18 3 31 13.5563 $w=2.02e-08 $l=2.3e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4860 $Y=0.0635 $X2=0.4860 $Y2=0.0405
r19 15 28 1.37684 $w=2.03185e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5125 $Y=0.0820 $X2=0.4990 $Y2=0.0820
r20 27 28 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.0820 $X2=0.4990 $Y2=0.0820
r21 27 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0820
+ $X2=0.4860 $Y2=0.0820
r22 26 27 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4750
+ $Y=0.0820 $X2=0.4860 $Y2=0.0820
r23 25 26 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4600
+ $Y=0.0820 $X2=0.4750 $Y2=0.0820
r24 24 25 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4310
+ $Y=0.0820 $X2=0.4600 $Y2=0.0820
r25 23 24 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.4145
+ $Y=0.0820 $X2=0.4310 $Y2=0.0820
r26 21 23 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4055
+ $Y=0.0820 $X2=0.4145 $Y2=0.0820
r27 12 21 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3965
+ $Y=0.0820 $X2=0.4055 $Y2=0.0820
r28 18 20 2.94116 $w=2.133e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.4060
+ $Y=0.0820 $X2=0.4160 $Y2=0.0820
r29 18 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4060 $Y=0.0820
+ $X2=0.4055 $Y2=0.0820
r30 1 18 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.3960
+ $Y=0.0820 $X2=0.4060 $Y2=0.0820
r31 1 19 0.851883 $w=1.865e-08 $l=2e-09 $layer=LIG $thickness=4.8e-08 $X=0.3960
+ $Y=0.0820 $X2=0.3940 $Y2=0.0820
r32 17 18 2.35044 $w=2.2e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.4050
+ $Y=0.0820 $X2=0.4060 $Y2=0.0820
r33 17 19 0.590723 $w=1.53e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4050 $Y=0.0820 $X2=0.3940 $Y2=0.0820
r34 17 20 0.590723 $w=1.53e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4050 $Y=0.0820 $X2=0.4160 $Y2=0.0820
r35 9 17 0.314665 $w=2.27e-07 $l=5.3e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4050 $Y2=0.0820
.ends

.subckt PM_ICGx1_ASAP7_75t_R%PD2 VSS 7 13 5 4 1
c1 1 VSS 0.00729323f
c2 4 VSS 0.00188005f
c3 5 VSS 0.00238554f
r1 13 12 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r2 5 12 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3800 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r3 10 5 9.87715 $w=2.32e-08 $l=2.1e-08 $layer=LISD $thickness=2.7e-08 $X=0.3570
+ $Y=0.2295 $X2=0.3780 $Y2=0.2295
r4 9 10 6.11443 $w=2.32e-08 $l=1.3e-08 $layer=LISD $thickness=2.7e-08 $X=0.3440
+ $Y=0.2295 $X2=0.3570 $Y2=0.2295
r5 8 9 2.82204 $w=2.32e-08 $l=6e-09 $layer=LISD $thickness=2.7e-08 $X=0.3380
+ $Y=0.2295 $X2=0.3440 $Y2=0.2295
r6 1 8 6.58477 $w=2.32e-08 $l=1.4e-08 $layer=LISD $thickness=2.7e-08 $X=0.3240
+ $Y=0.2295 $X2=0.3380 $Y2=0.2295
r7 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2295 $X2=0.3220 $Y2=0.2295
r8 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2295 $X2=0.3095 $Y2=0.2295
.ends

.subckt PM_ICGx1_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.00364748f
.ends

.subckt PM_ICGx1_ASAP7_75t_R%GCLKN VSS 12 40 41 49 50 53 54 13 14 3 16 5 4 15
+ 17 20 1 19 22 21
c1 1 VSS 0.00372511f
c2 3 VSS 0.00842433f
c3 4 VSS 0.00519575f
c4 5 VSS 0.00816282f
c5 12 VSS 0.0795253f
c6 13 VSS 0.00294664f
c7 14 VSS 0.00393829f
c8 15 VSS 0.00393305f
c9 16 VSS 0.0122393f
c10 17 VSS 0.00584557f
c11 18 VSS 0.00137576f
c12 19 VSS 0.00162224f
c13 20 VSS 0.00352744f
c14 21 VSS 0.000497481f
c15 22 VSS 0.00059592f
r1 54 52 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.2160 $X2=0.7165 $Y2=0.2160
r2 3 52 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7020 $Y=0.2160 $X2=0.7165 $Y2=0.2160
r3 14 3 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.2160 $X2=0.7020 $Y2=0.2160
r4 53 14 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.2160 $X2=0.6875 $Y2=0.2160
r5 50 48 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8270 $Y=0.2160 $X2=0.8245 $Y2=0.2160
r6 5 48 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8100 $Y=0.2160 $X2=0.8245 $Y2=0.2160
r7 15 5 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.2160 $X2=0.8100 $Y2=0.2160
r8 49 15 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.2160 $X2=0.7955 $Y2=0.2160
r9 3 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7020 $Y=0.2160
+ $X2=0.7020 $Y2=0.2310
r10 5 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8100 $Y=0.2160
+ $X2=0.8100 $Y2=0.2310
r11 45 46 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.2310 $X2=0.7380 $Y2=0.2310
r12 42 43 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.2310 $X2=0.8235 $Y2=0.2310
r13 16 42 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.2310 $X2=0.8100 $Y2=0.2310
r14 16 46 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.2310 $X2=0.7380 $Y2=0.2310
r15 40 39 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.0675 $X2=0.7705 $Y2=0.0675
r16 4 39 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7560 $Y=0.0675 $X2=0.7705 $Y2=0.0675
r17 13 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7415 $Y=0.0675 $X2=0.7560 $Y2=0.0675
r18 41 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.0675 $X2=0.7415 $Y2=0.0675
r19 36 43 1.20242 $w=1.425e-08 $l=1.54434e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8370 $Y=0.2235 $X2=0.8235 $Y2=0.2310
r20 35 36 2.01858 $w=1.37895e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.8370 $Y=0.2140 $X2=0.8370 $Y2=0.2235
r21 34 35 2.37574 $w=1.49231e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8370 $Y=0.2010 $X2=0.8370 $Y2=0.2140
r22 20 34 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1920 $X2=0.8370 $Y2=0.2010
r23 4 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7560 $Y=0.0675
+ $X2=0.7560 $Y2=0.0720
r24 18 22 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8640 $Y=0.1970 $X2=0.8910 $Y2=0.1970
r25 18 20 4.60559 $w=1.39091e-08 $l=2.74591e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8640 $Y=0.1970 $X2=0.8370 $Y2=0.1920
r26 32 33 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.0720 $X2=0.7965 $Y2=0.0720
r27 30 33 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.0720 $X2=0.7965 $Y2=0.0720
r28 29 30 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.8625
+ $Y=0.0720 $X2=0.8370 $Y2=0.0720
r29 17 21 0.79938 $w=1.72857e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8805 $Y=0.0720 $X2=0.8910 $Y2=0.0720
r30 17 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8805
+ $Y=0.0720 $X2=0.8625 $Y2=0.0720
r31 22 28 5.22999 $w=1.59898e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8910 $Y=0.1970 $X2=0.8910 $Y2=0.1675
r32 21 27 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.0720 $X2=0.8910 $Y2=0.0900
r33 26 28 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1460 $X2=0.8910 $Y2=0.1675
r34 25 26 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1360 $X2=0.8910 $Y2=0.1460
r35 19 25 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1130 $X2=0.8910 $Y2=0.1360
r36 19 27 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1130 $X2=0.8910 $Y2=0.0900
r37 12 1 6.51726 $w=1.18568e-07 $l=5e-10 $layer=LIG $thickness=5.19024e-08
+ $X=0.8910 $Y=0.1350 $X2=0.8910 $Y2=0.1355
r38 1 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8910 $Y=0.1355
+ $X2=0.8910 $Y2=0.1360
.ends

.subckt PM_ICGx1_ASAP7_75t_R%CLKN VSS 9 51 53 10 17 12 3 14 1 13 11 16 15 4
c1 1 VSS 0.000109604f
c2 3 VSS 0.00618368f
c3 4 VSS 0.00786232f
c4 9 VSS 0.00447113f
c5 10 VSS 0.00596062f
c6 11 VSS 0.00598824f
c7 12 VSS 0.00182112f
c8 13 VSS 0.00120214f
c9 14 VSS 0.000631452f
c10 15 VSS 0.000854063f
c11 16 VSS 0.00629182f
c12 17 VSS 0.00866892f
r1 53 52 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.2025 $X2=0.6085 $Y2=0.2025
r2 11 52 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5960 $Y=0.2025 $X2=0.6085 $Y2=0.2025
r3 51 50 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.0675 $X2=0.6085 $Y2=0.0675
r4 10 50 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5960 $Y=0.0675 $X2=0.6085 $Y2=0.0675
r5 4 44 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2295
+ $X2=0.5940 $Y2=0.2320
r6 3 41 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0605
+ $X2=0.5940 $Y2=0.0860
r7 43 44 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5810
+ $Y=0.2320 $X2=0.5940 $Y2=0.2320
r8 16 39 1.03499 $w=1.77368e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.5680 $Y=0.2320 $X2=0.5680 $Y2=0.2225
r9 16 43 1.85116 $w=1.64615e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5680 $Y=0.2320 $X2=0.5810 $Y2=0.2320
r10 40 41 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5810
+ $Y=0.0860 $X2=0.5940 $Y2=0.0860
r11 15 36 3.36689 $w=1.53077e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5680 $Y=0.0860 $X2=0.5680 $Y2=0.1055
r12 15 40 1.85116 $w=1.64615e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5680 $Y=0.0860 $X2=0.5810 $Y2=0.0860
r13 38 39 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5680
+ $Y=0.2100 $X2=0.5680 $Y2=0.2225
r14 37 38 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5680
+ $Y=0.1970 $X2=0.5680 $Y2=0.2100
r15 35 37 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5680
+ $Y=0.1880 $X2=0.5680 $Y2=0.1970
r16 13 35 9.32759 $w=1.3e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.5680
+ $Y=0.1480 $X2=0.5680 $Y2=0.1880
r17 13 36 9.91056 $w=1.3e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5680
+ $Y=0.1480 $X2=0.5680 $Y2=0.1055
r18 33 35 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.5680 $Y=0.1890
+ $X2=0.5680 $Y2=0.1880
r19 32 33 30.0815 $w=1.3e-08 $l=1.29e-07 $layer=M2 $thickness=3.6e-08 $X=0.4390
+ $Y=0.1890 $X2=0.5680 $Y2=0.1890
r20 31 32 30.0815 $w=1.3e-08 $l=1.29e-07 $layer=M2 $thickness=3.6e-08 $X=0.3100
+ $Y=0.1890 $X2=0.4390 $Y2=0.1890
r21 17 31 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.2985
+ $Y=0.1890 $X2=0.3100 $Y2=0.1890
r22 29 31 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.3145 $Y=0.1890
+ $X2=0.3100 $Y2=0.1890
r23 28 29 1.51573 $w=1.3e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3080
+ $Y=0.1890 $X2=0.3145 $Y2=0.1890
r24 27 28 0.721491 $w=1.57778e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.3035 $Y=0.1890 $X2=0.3080 $Y2=0.1890
r25 14 27 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2945
+ $Y=0.1890 $X2=0.3035 $Y2=0.1890
r26 26 27 4.68572 $w=1.35814e-08 $l=2.87446e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1610 $X2=0.3035 $Y2=0.1890
r27 25 26 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1330 $X2=0.2970 $Y2=0.1610
r28 24 25 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1215 $X2=0.2970 $Y2=0.1330
r29 12 24 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0955 $X2=0.2970 $Y2=0.1215
r30 1 21 2.88023 $w=2.1e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.2970
+ $Y=0.1335 $X2=0.2970 $Y2=0.1335
r31 1 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1335
+ $X2=0.2970 $Y2=0.1330
r32 9 21 0.314665 $w=2.27e-07 $l=1.5e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2970 $Y2=0.1335
r33 4 11 1e-05
r34 3 10 1e-05
.ends

.subckt PM_ICGx1_ASAP7_75t_R%CLK VSS 54 10 11 12 13 14 23 1 15 21 20 16 8 17 3
+ 2 19 22 4 18
c1 1 VSS 0.00397182f
c2 2 VSS 0.00191704f
c3 3 VSS 0.00748125f
c4 4 VSS 0.00902009f
c5 8 VSS 0.00410516f
c6 10 VSS 0.00633535f
c7 11 VSS 0.0063201f
c8 12 VSS 0.0821357f
c9 13 VSS 0.0342954f
c10 14 VSS 0.0343942f
c11 15 VSS 0.00485748f
c12 16 VSS 0.00472506f
c13 17 VSS 0.00493357f
c14 18 VSS 0.00230895f
c15 19 VSS 0.00200773f
c16 20 VSS 0.00396944f
c17 21 VSS 0.00251798f
c18 22 VSS 0.00247764f
c19 23 VSS 0.00599892f
r1 2 78 3.16825 $w=2.1e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.3520
+ $Y=0.1335 $X2=0.3555 $Y2=0.1335
r2 11 2 3.48292 $w=1.19095e-07 $l=1.80278e-09 $layer=LIG $thickness=5.18095e-08
+ $X=0.3510 $Y=0.1350 $X2=0.3520 $Y2=0.1335
r3 77 78 4.91375 $w=2.12e-08 $l=1.5e-09 $layer=LISD $thickness=2.7e-08
+ $X=0.3570 $Y=0.1335 $X2=0.3555 $Y2=0.1335
r4 76 77 11.4654 $w=2.12e-08 $l=2.1e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.3780 $Y=0.1335 $X2=0.3570 $Y2=0.1335
r5 75 76 7.37062 $w=2.12e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.3915 $Y=0.1335 $X2=0.3780 $Y2=0.1335
r6 8 73 5.7327 $w=2.12e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08 $X=0.3945
+ $Y=0.1335 $X2=0.4050 $Y2=0.1335
r7 8 75 1.63792 $w=2.12e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.3945
+ $Y=0.1335 $X2=0.3915 $Y2=0.1335
r8 1 62 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1335
+ $X2=0.2430 $Y2=0.1330
r9 10 1 3.19489 $w=1.24e-07 $l=1.5e-09 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1335
r10 69 70 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1340 $X2=0.4050 $Y2=0.1435
r11 69 73 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4050 $Y=0.1340
+ $X2=0.4050 $Y2=0.1335
r12 19 20 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1530 $X2=0.4230 $Y2=0.1530
r13 19 70 1.03499 $w=1.77368e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.1530 $X2=0.4050 $Y2=0.1435
r14 63 64 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1430 $X2=0.2430 $Y2=0.1530
r15 62 63 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1330 $X2=0.2430 $Y2=0.1430
r16 15 62 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1215 $X2=0.2430 $Y2=0.1330
r17 20 52 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4230 $Y=0.1530
+ $X2=0.4230 $Y2=0.1530
r18 3 46 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6210 $Y=0.1350
+ $X2=0.6210 $Y2=0.1330
r19 12 3 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1350
r20 57 58 7.22888 $w=1.3e-08 $l=3.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1530 $X2=0.2740 $Y2=0.1530
r21 57 64 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.2430 $Y=0.1530
+ $X2=0.2430 $Y2=0.1530
r22 54 55 1.10765 $w=1.3e-08 $l=4.7e-09 $layer=M2 $thickness=3.6e-08 $X=0.5730
+ $Y=0.1530 $X2=0.5777 $Y2=0.1530
r23 54 53 16.4982 $w=1.3e-08 $l=7.08e-08 $layer=M2 $thickness=3.6e-08 $X=0.5730
+ $Y=0.1530 $X2=0.5022 $Y2=0.1530
r24 52 53 18.4803 $w=1.3e-08 $l=7.92e-08 $layer=M2 $thickness=3.6e-08 $X=0.4230
+ $Y=0.1530 $X2=0.5022 $Y2=0.1530
r25 51 52 15.8569 $w=1.3e-08 $l=6.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.3550
+ $Y=0.1530 $X2=0.4230 $Y2=0.1530
r26 51 58 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.3550
+ $Y=0.1530 $X2=0.2740 $Y2=0.1530
r27 23 49 5.59655 $w=1.3e-08 $l=2.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.5970
+ $Y=0.1530 $X2=0.6210 $Y2=0.1530
r28 23 55 4.4889 $w=1.3e-08 $l=1.93e-08 $layer=M2 $thickness=3.6e-08 $X=0.5970
+ $Y=0.1530 $X2=0.5777 $Y2=0.1530
r29 47 48 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1430 $X2=0.6210 $Y2=0.1455
r30 46 47 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1330 $X2=0.6210 $Y2=0.1430
r31 16 44 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1545 $X2=0.6210 $Y2=0.1700
r32 16 48 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1545 $X2=0.6210 $Y2=0.1455
r33 16 49 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.6210 $Y=0.1545
+ $X2=0.6210 $Y2=0.1530
r34 21 43 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.1870 $X2=0.6480 $Y2=0.1870
r35 21 44 2.31511 $w=1.81882e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.1870 $X2=0.6210 $Y2=0.1700
r36 42 43 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1870 $X2=0.6480 $Y2=0.1870
r37 41 42 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6860
+ $Y=0.1870 $X2=0.6750 $Y2=0.1870
r38 17 22 7.38932 $w=1.37246e-08 $l=3.87072e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7175 $Y=0.1870 $X2=0.7560 $Y2=0.1830
r39 17 41 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.7175
+ $Y=0.1870 $X2=0.6860 $Y2=0.1870
r40 22 38 1.32639 $w=1.59412e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.7560 $Y=0.1830 $X2=0.7560 $Y2=0.1745
r41 13 33 2.92627 $w=1.245e-07 $l=2.7e-08 $layer=LIG $thickness=5.2e-08
+ $X=0.7290 $Y=0.1350 $X2=0.7290 $Y2=0.1620
r42 37 38 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.1620 $X2=0.7560 $Y2=0.1745
r43 36 37 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.1500 $X2=0.7560 $Y2=0.1620
r44 18 36 1.28254 $w=1.3e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.1445 $X2=0.7560 $Y2=0.1500
r45 31 33 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7415 $Y=0.1620 $X2=0.7290 $Y2=0.1620
r46 30 31 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7560 $Y=0.1620 $X2=0.7415 $Y2=0.1620
r47 30 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7560 $Y=0.1620
+ $X2=0.7560 $Y2=0.1620
r48 29 30 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7705 $Y=0.1620 $X2=0.7560 $Y2=0.1620
r49 4 28 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.7830
+ $Y=0.1620 $X2=0.7830 $Y2=0.1620
r50 4 29 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7830 $Y=0.1620 $X2=0.7705 $Y2=0.1620
r51 4 35 2.90696 $w=2.1681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7830 $Y=0.1620 $X2=0.7935 $Y2=0.1620
r52 28 29 1.47681 $w=1.53e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7830 $Y=0.1620 $X2=0.7705 $Y2=0.1620
r53 28 35 0.295362 $w=1.53e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7830 $Y=0.1620 $X2=0.7935 $Y2=0.1620
r54 14 28 0.314665 $w=2.27e-07 $l=2.7e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.7830 $Y=0.1350 $X2=0.7830 $Y2=0.1620
.ends

.subckt PM_ICGx1_ASAP7_75t_R%MH VSS 13 14 15 76 80 98 102 23 21 7 19 29 17 27
+ 32 33 18 3 1 25 26 20 22 24 16 8 2 30 31
c1 1 VSS 0.0023512f
c2 2 VSS 0.0046007f
c3 3 VSS 0.00407688f
c4 7 VSS 0.00514597f
c5 8 VSS 0.00508077f
c6 13 VSS 0.036861f
c7 14 VSS 0.0818819f
c8 15 VSS 0.081877f
c9 16 VSS 0.00317768f
c10 17 VSS 0.000556973f
c11 18 VSS 0.00315418f
c12 19 VSS 0.000592325f
c13 20 VSS 0.00829057f
c14 21 VSS 0.00384165f
c15 22 VSS 0.000842461f
c16 23 VSS 0.00042682f
c17 24 VSS 0.0293067f
c18 25 VSS 0.00200943f
c19 26 VSS 0.00222539f
c20 27 VSS 0.00204787f
c21 28 VSS 0.00225312f
c22 29 VSS 7.69109e-20
c23 30 VSS 0.00263409f
c24 31 VSS 0.00334412f
c25 32 VSS 0.000693341f
c26 33 VSS 0.00136101f
r1 102 101 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2295 $X2=0.2845 $Y2=0.2295
r2 100 101 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2800 $Y=0.2295 $X2=0.2845 $Y2=0.2295
r3 18 100 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2680 $Y=0.2295 $X2=0.2800 $Y2=0.2295
r4 19 18 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2295 $X2=0.2680 $Y2=0.2295
r5 96 97 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.1890 $X2=0.2600 $Y2=0.1890
r6 98 96 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.1890 $X2=0.2555 $Y2=0.1890
r7 18 97 0.185185 $w=5.4e-08 $l=1e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.1890 $X2=0.2600 $Y2=0.1890
r8 7 93 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2295
+ $X2=0.2700 $Y2=0.2320
r9 7 18 23.8708 $w=2.02e-08 $l=4.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.2700 $Y=0.2295 $X2=0.2700 $Y2=0.1890
r10 93 94 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2320 $X2=0.2835 $Y2=0.2320
r11 91 94 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3060
+ $Y=0.2320 $X2=0.2835 $Y2=0.2320
r12 20 30 2.96589 $w=1.31923e-08 $l=2.31193e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3365 $Y=0.2320 $X2=0.3580 $Y2=0.2235
r13 20 91 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.3365
+ $Y=0.2320 $X2=0.3060 $Y2=0.2320
r14 1 85 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1900
+ $X2=0.4590 $Y2=0.1900
r15 13 1 3.49039 $w=1.235e-07 $l=5.5e-08 $layer=LIG $thickness=5.2e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4590 $Y2=0.1900
r16 23 74 2.8493 $w=1.32e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.2110 $X2=0.3580 $Y2=0.1985
r17 23 30 2.8493 $w=1.32e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.2110 $X2=0.3580 $Y2=0.2235
r18 84 85 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4485
+ $Y=0.1900 $X2=0.4590 $Y2=0.1900
r19 83 84 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4305
+ $Y=0.1900 $X2=0.4485 $Y2=0.1900
r20 82 83 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1900 $X2=0.4305 $Y2=0.1900
r21 81 82 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3940
+ $Y=0.1900 $X2=0.4050 $Y2=0.1900
r22 25 29 3.78225 $w=1.50238e-08 $l=2.15058e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3795 $Y=0.1900 $X2=0.3580 $Y2=0.1895
r23 25 81 3.38125 $w=1.3e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3795
+ $Y=0.1900 $X2=0.3940 $Y2=0.1900
r24 80 79 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0405 $X2=0.3385 $Y2=0.0405
r25 78 79 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3340 $Y=0.0405 $X2=0.3385 $Y2=0.0405
r26 8 78 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3220 $Y=0.0405 $X2=0.3340 $Y2=0.0405
r27 17 8 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0405 $X2=0.3220 $Y2=0.0405
r28 16 8 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0810 $X2=0.3220 $Y2=0.0810
r29 76 16 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0810 $X2=0.3095 $Y2=0.0810
r30 29 69 0.983973 $w=1.77222e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.3580 $Y=0.1895 $X2=0.3580 $Y2=0.1805
r31 29 74 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.1895 $X2=0.3580 $Y2=0.1985
r32 8 63 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0405
+ $X2=0.3195 $Y2=0.0360
r33 68 69 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.1710 $X2=0.3580 $Y2=0.1805
r34 67 68 6.99569 $w=1.3e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.1410 $X2=0.3580 $Y2=0.1710
r35 66 67 8.27824 $w=1.3e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.1055 $X2=0.3580 $Y2=0.1410
r36 65 66 5.47996 $w=1.3e-08 $l=2.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.0820 $X2=0.3580 $Y2=0.1055
r37 64 65 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.0725 $X2=0.3580 $Y2=0.0820
r38 22 28 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.0585 $X2=0.3580 $Y2=0.0360
r39 22 64 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.0585 $X2=0.3580 $Y2=0.0725
r40 21 61 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3285
+ $Y=0.0360 $X2=0.3410 $Y2=0.0360
r41 21 63 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3285
+ $Y=0.0360 $X2=0.3195 $Y2=0.0360
r42 28 60 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3580 $Y=0.0360 $X2=0.3795 $Y2=0.0360
r43 28 61 2.78392 $w=1.56471e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3580 $Y=0.0360 $X2=0.3410 $Y2=0.0360
r44 59 60 18.0722 $w=1.3e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.4570
+ $Y=0.0360 $X2=0.3795 $Y2=0.0360
r45 58 59 19.4713 $w=1.3e-08 $l=8.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5405
+ $Y=0.0360 $X2=0.4570 $Y2=0.0360
r46 57 58 10.1438 $w=1.3e-08 $l=4.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5840
+ $Y=0.0360 $X2=0.5405 $Y2=0.0360
r47 56 57 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.6105
+ $Y=0.0360 $X2=0.5840 $Y2=0.0360
r48 55 56 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0360 $X2=0.6105 $Y2=0.0360
r49 24 31 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6480 $Y=0.0360 $X2=0.6750 $Y2=0.0360
r50 24 55 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.6480
+ $Y=0.0360 $X2=0.6210 $Y2=0.0360
r51 31 51 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0360 $X2=0.6750 $Y2=0.0540
r52 2 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6750 $Y=0.1350
+ $X2=0.6750 $Y2=0.1330
r53 14 2 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6750
+ $Y=0.1350 $X2=0.6750 $Y2=0.1350
r54 50 51 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0680 $X2=0.6750 $Y2=0.0540
r55 49 50 1.63233 $w=1.3e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0750 $X2=0.6750 $Y2=0.0680
r56 48 49 0.932759 $w=1.3e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0790 $X2=0.6750 $Y2=0.0750
r57 47 48 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0880 $X2=0.6750 $Y2=0.0790
r58 26 32 1.33376 $w=1.70476e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6750 $Y=0.0970 $X2=0.6750 $Y2=0.1075
r59 26 47 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0970 $X2=0.6750 $Y2=0.0880
r60 44 45 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1205 $X2=0.6750 $Y2=0.1330
r61 43 44 0.867186 $w=1.3625e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.6750 $Y=0.1165 $X2=0.6750 $Y2=0.1205
r62 32 43 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1075 $X2=0.6750 $Y2=0.1165
r63 42 43 6.81353 $w=1.30847e-08 $l=3.89391e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7130 $Y=0.1080 $X2=0.6750 $Y2=0.1165
r64 41 42 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.7445
+ $Y=0.1080 $X2=0.7130 $Y2=0.1080
r65 40 41 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.1080 $X2=0.7445 $Y2=0.1080
r66 27 38 8.26388 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7965 $Y=0.1080 $X2=0.8370 $Y2=0.1080
r67 27 40 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.7965
+ $Y=0.1080 $X2=0.7560 $Y2=0.1080
r68 33 37 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1205 $X2=0.8370 $Y2=0.1330
r69 33 38 1.73456 $w=1.66e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8370 $Y=0.1205 $X2=0.8370 $Y2=0.1080
r70 15 3 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.8370
+ $Y=0.1350 $X2=0.8370 $Y2=0.1350
r71 3 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8370 $Y=0.1350
+ $X2=0.8370 $Y2=0.1330
.ends


*
.SUBCKT ICGx1_ASAP7_75t_R VSS VDD ENA SE CLK GCLK
*
* VSS VSS
* VDD VDD
* ENA ENA
* SE SE
* CLK CLK
* GCLK GCLK
*
*

MM19 N_MM19_d N_MM19_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM27 N_MM27_d N_MM18_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM10_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM6 N_MM6_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM20 N_MM20_d N_MM21_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM14 N_MM14_d N_MM0_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM16_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM13 N_MM13_d N_MM13_g N_MM13_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM12 N_MM12_d N_MM12_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24 N_MM24_d N_MM24_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM26 N_MM26_d N_MM19_g N_MM26_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM18 N_MM18_d N_MM18_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM21 N_MM21_d N_MM21_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM16 N_MM16_d N_MM16_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM16@2 N_MM16@2_d N_MM13_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM0@2 N_MM0@2_d N_MM12_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM25 N_MM25_d N_MM24_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "ICGx1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "ICGx1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_ICGx1_ASAP7_75t_R%NOS1 VSS N_MM26_s N_MM18_d N_NOS1_1
+ PM_ICGx1_ASAP7_75t_R%NOS1
cc_1 N_NOS1_1 N_MM19_g 0.0125299f
cc_2 N_NOS1_1 N_MM18_g 0.0125764f
x_PM_ICGx1_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_ICGx1_ASAP7_75t_R%noxref_20
cc_3 N_noxref_20_1 N_MM19_g 0.00393299f
cc_4 N_noxref_20_1 N_NET0121_11 0.0276625f
cc_5 N_noxref_20_1 N_noxref_19_1 0.00208912f
x_PM_ICGx1_ASAP7_75t_R%SE VSS SE N_MM18_g N_SE_1 N_SE_4 PM_ICGx1_ASAP7_75t_R%SE
cc_6 N_SE_1 N_ENA_1 0.001696f
cc_7 N_SE_4 N_ENA_4 0.00520432f
cc_8 N_MM18_g N_MM19_g 0.00985303f
x_PM_ICGx1_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_ICGx1_ASAP7_75t_R%noxref_19
cc_9 N_noxref_19_1 N_MM19_g 0.00394103f
cc_10 N_noxref_19_1 N_NET0121_10 0.000403813f
x_PM_ICGx1_ASAP7_75t_R%ENA VSS ENA N_MM19_g N_ENA_1 N_ENA_4
+ PM_ICGx1_ASAP7_75t_R%ENA
x_PM_ICGx1_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_ICGx1_ASAP7_75t_R%noxref_25
cc_11 N_noxref_25_1 N_MM24_g 0.00145656f
cc_12 N_noxref_25_1 N_GCLK_7 0.0386109f
x_PM_ICGx1_ASAP7_75t_R%noxref_26 VSS N_noxref_26_1
+ PM_ICGx1_ASAP7_75t_R%noxref_26
cc_13 N_noxref_26_1 N_MM24_g 0.00145336f
cc_14 N_noxref_26_1 N_GCLK_8 0.0384583f
cc_15 N_noxref_26_1 N_noxref_25_1 0.00177505f
x_PM_ICGx1_ASAP7_75t_R%GCLK VSS GCLK N_MM24_d N_MM25_d N_GCLK_7 N_GCLK_9
+ N_GCLK_1 N_GCLK_2 N_GCLK_8 N_GCLK_10 N_GCLK_11 PM_ICGx1_ASAP7_75t_R%GCLK
cc_16 N_GCLK_7 N_GCLKN_1 0.000786068f
cc_17 N_GCLK_9 N_GCLKN_17 0.000874322f
cc_18 N_GCLK_1 N_MM24_g 0.00142726f
cc_19 N_GCLK_2 N_MM24_g 0.00145604f
cc_20 N_GCLK_8 N_GCLKN_1 0.00179436f
cc_21 N_GCLK_10 N_GCLKN_22 0.00226495f
cc_22 N_GCLK_9 N_GCLKN_21 0.00288808f
cc_23 N_GCLK_8 N_MM24_g 0.0151737f
cc_24 N_GCLK_11 N_GCLKN_19 0.00596823f
cc_25 N_GCLK_7 N_MM24_g 0.0554376f
x_PM_ICGx1_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_ICGx1_ASAP7_75t_R%noxref_24
cc_26 N_noxref_24_1 N_MM21_g 0.00136833f
cc_27 N_noxref_24_1 N_CLKN_4 0.00041051f
cc_28 N_noxref_24_1 N_CLKN_11 0.0373745f
cc_29 N_noxref_24_1 N_MS_11 0.000538342f
cc_30 N_noxref_24_1 N_noxref_21_1 0.000473222f
cc_31 N_noxref_24_1 N_noxref_22_1 0.00777072f
cc_32 N_noxref_24_1 N_noxref_23_1 0.0012309f
x_PM_ICGx1_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_ICGx1_ASAP7_75t_R%noxref_23
cc_33 N_noxref_23_1 N_MM21_g 0.0013639f
cc_34 N_noxref_23_1 N_CLKN_10 0.0376345f
cc_35 N_noxref_23_1 N_MS_10 0.000574231f
cc_36 N_noxref_23_1 N_noxref_21_1 0.00772764f
cc_37 N_noxref_23_1 N_noxref_22_1 0.000477044f
x_PM_ICGx1_ASAP7_75t_R%NET0121 VSS N_MM3_g N_MM19_d N_MM27_d N_MM26_d
+ N_NET0121_11 N_NET0121_13 N_NET0121_4 N_NET0121_3 N_NET0121_12 N_NET0121_10
+ N_NET0121_1 N_NET0121_14 PM_ICGx1_ASAP7_75t_R%NET0121
cc_38 N_NET0121_11 N_ENA_1 0.000579346f
cc_39 N_NET0121_13 N_ENA_4 0.000725209f
cc_40 N_NET0121_4 N_MM19_g 0.000750771f
cc_41 N_NET0121_3 N_MM19_g 0.00108943f
cc_42 N_NET0121_12 N_ENA_4 0.00143521f
cc_43 N_NET0121_4 N_ENA_4 0.00304002f
cc_44 N_NET0121_11 N_MM19_g 0.0111053f
cc_45 N_NET0121_10 N_MM19_g 0.0403174f
cc_46 N_NET0121_1 N_MM18_g 0.000968072f
cc_47 N_NET0121_13 N_SE_4 0.00103806f
cc_48 N_NET0121_1 N_SE_1 0.00119164f
cc_49 N_NET0121_12 N_SE_4 0.00121383f
cc_50 N_NET0121_10 N_MM18_g 0.0109236f
cc_51 N_NET0121_14 N_SE_4 0.00764419f
cc_52 N_MM3_g N_MM18_g 0.0186741f
x_PM_ICGx1_ASAP7_75t_R%PD1 VSS N_MM5_d N_MM4_s N_PD1_4 N_PD1_5 N_PD1_1
+ PM_ICGx1_ASAP7_75t_R%PD1
cc_53 N_PD1_4 N_NET0121_14 0.000812593f
cc_54 N_PD1_4 N_MM3_g 0.0359859f
cc_55 N_PD1_5 N_CLK_1 0.00236641f
cc_56 N_PD1_5 N_MM1_g 0.0731249f
cc_57 N_PD1_5 N_CLKN_12 0.000624267f
cc_58 N_PD1_5 N_CLKN_1 0.00068583f
cc_59 N_PD1_5 N_MM10_g 0.0346182f
cc_60 N_PD1_1 N_MH_8 0.00134665f
cc_61 N_PD1_1 N_MH_16 0.00300365f
x_PM_ICGx1_ASAP7_75t_R%NET0140 VSS N_MM14_d N_MM2_s N_NET0140_1
+ PM_ICGx1_ASAP7_75t_R%NET0140
cc_62 N_NET0140_1 N_MM16_g 0.0174401f
cc_63 N_NET0140_1 N_MM0_g 0.017269f
x_PM_ICGx1_ASAP7_75t_R%PU1 VSS N_MM3_d N_MM1_s N_PU1_3 N_PU1_1
+ PM_ICGx1_ASAP7_75t_R%PU1
cc_64 N_PU1_3 N_NET0121_1 0.000627883f
cc_65 N_PU1_3 N_MM3_g 0.0348942f
cc_66 N_PU1_3 N_CLK_15 0.000339666f
cc_67 N_PU1_3 N_CLK_1 0.000513615f
cc_68 N_PU1_3 N_MM1_g 0.0336019f
cc_69 N_PU1_1 N_MH_18 0.00109742f
cc_70 N_PU1_1 N_MH_7 0.00288867f
x_PM_ICGx1_ASAP7_75t_R%PD3 VSS N_MM9_s N_MM8_d N_PD3_3 N_PD3_1
+ PM_ICGx1_ASAP7_75t_R%PD3
cc_71 N_PD3_3 N_MM9_g 0.0146829f
cc_72 N_PD3_3 N_MM11_g 0.0162452f
cc_73 N_PD3_1 N_MH_22 0.00019306f
cc_74 N_PD3_1 N_MH_16 0.000612332f
cc_75 N_PD3_1 N_MH_24 0.000308143f
cc_76 N_PD3_1 N_MH_8 0.00210846f
x_PM_ICGx1_ASAP7_75t_R%NET0141 VSS N_MM13_s N_MM12_d N_NET0141_1
+ PM_ICGx1_ASAP7_75t_R%NET0141
cc_77 N_NET0141_1 N_MM13_g 0.0173257f
cc_78 N_NET0141_1 N_MM12_g 0.0173386f
x_PM_ICGx1_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_ICGx1_ASAP7_75t_R%noxref_21
cc_79 N_noxref_21_1 N_CLKN_10 0.000837518f
cc_80 N_noxref_21_1 N_MS_3 0.00100914f
cc_81 N_noxref_21_1 N_MS_10 0.0169534f
cc_82 N_noxref_21_1 N_MM7_g 0.00534817f
x_PM_ICGx1_ASAP7_75t_R%MS VSS N_MM11_g N_MM6_d N_MM7_d N_MS_1 N_MS_12 N_MS_13
+ N_MS_15 N_MS_3 N_MS_14 N_MS_4 N_MS_11 N_MS_10 PM_ICGx1_ASAP7_75t_R%MS
cc_83 N_MM11_g N_CLK_20 0.000217534f
cc_84 N_MM11_g N_CLK_23 0.000125382f
cc_85 N_MM11_g N_CLK_8 0.00293903f
cc_86 N_MS_1 N_CLK_19 0.000552116f
cc_87 N_MS_1 N_CLK_8 0.00153715f
cc_88 N_MS_12 N_CLK_20 0.000626225f
cc_89 N_MS_13 N_CLK_23 0.00150957f
cc_90 N_MS_12 N_CLK_23 0.0016024f
cc_91 N_MS_12 N_CLK_19 0.00255848f
cc_92 N_MM11_g N_MM9_g 0.013171f
cc_93 N_MS_13 N_CLKN_11 0.000122571f
cc_94 N_MS_13 N_CLKN_15 0.000221069f
cc_95 N_MS_15 N_CLKN_3 0.00024744f
cc_96 N_MS_3 N_CLKN_15 0.000253119f
cc_97 N_MS_13 N_CLKN_4 0.000275436f
cc_98 N_MS_14 N_CLKN_16 0.000855618f
cc_99 N_MS_15 N_CLKN_15 0.000951897f
cc_100 N_MS_14 N_CLKN_17 0.00148256f
cc_101 N_MS_13 N_CLKN_13 0.00668115f
x_PM_ICGx1_ASAP7_75t_R%PD2 VSS N_MM10_s N_MM11_d N_PD2_5 N_PD2_4 N_PD2_1
+ PM_ICGx1_ASAP7_75t_R%PD2
cc_102 N_PD2_5 N_CLK_8 0.000221014f
cc_103 N_PD2_4 N_MM9_g 0.00732318f
cc_104 N_PD2_1 N_MM9_g 0.000993918f
cc_105 N_PD2_5 N_MM9_g 0.023718f
cc_106 N_PD2_1 N_MM10_g 0.000492679f
cc_107 N_PD2_4 N_MM10_g 0.0149734f
cc_108 N_PD2_5 N_MM11_g 0.0149323f
cc_109 N_PD2_1 N_MH_29 0.00010106f
cc_110 N_PD2_1 N_MH_7 0.000117213f
cc_111 N_PD2_1 N_MH_23 0.000256157f
cc_112 N_PD2_1 N_MH_25 0.000296436f
cc_113 N_PD2_4 N_MH_18 0.000643057f
cc_114 N_PD2_1 N_MH_20 0.000491767f
cc_115 N_PD2_4 N_MH_7 0.000618656f
cc_116 N_PD2_1 N_MH_30 0.00270059f
x_PM_ICGx1_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_ICGx1_ASAP7_75t_R%noxref_22
cc_117 N_noxref_22_1 N_CLKN_11 0.000956656f
cc_118 N_noxref_22_1 N_MS_11 0.0170564f
cc_119 N_noxref_22_1 N_MM7_g 0.00577904f
cc_120 N_noxref_22_1 N_noxref_21_1 0.00153657f
x_PM_ICGx1_ASAP7_75t_R%GCLKN VSS N_MM24_g N_MM13_d N_MM2_d N_MM16@2_d N_MM0@2_d
+ N_MM0_d N_MM16_d N_GCLKN_13 N_GCLKN_14 N_GCLKN_3 N_GCLKN_16 N_GCLKN_5
+ N_GCLKN_4 N_GCLKN_15 N_GCLKN_17 N_GCLKN_20 N_GCLKN_1 N_GCLKN_19 N_GCLKN_22
+ N_GCLKN_21 PM_ICGx1_ASAP7_75t_R%GCLKN
cc_121 N_GCLKN_13 N_CLK_22 0.000397519f
cc_122 N_GCLKN_13 N_CLK_23 0.000171454f
cc_123 N_GCLKN_13 N_CLK_18 0.000289281f
cc_124 N_GCLKN_13 N_CLK_4 0.000339561f
cc_125 N_GCLKN_14 N_MM16_g 0.011491f
cc_126 N_GCLKN_3 N_CLK_17 0.000418501f
cc_127 N_GCLKN_16 N_CLK_18 0.00047467f
cc_128 N_GCLKN_5 N_MM13_g 0.000844971f
cc_129 N_GCLKN_3 N_MM16_g 0.00125952f
cc_130 N_GCLKN_4 N_MM13_g 0.00149906f
cc_131 N_GCLKN_15 N_CLK_4 0.00245486f
cc_132 N_GCLKN_16 N_CLK_17 0.00251809f
cc_133 N_GCLKN_16 N_CLK_22 0.0038446f
cc_134 N_GCLKN_15 N_MM13_g 0.0109476f
cc_135 N_GCLKN_13 N_MM16_g 0.0331132f
cc_136 N_GCLKN_13 N_MM13_g 0.0655197f
cc_137 N_GCLKN_14 N_MH_2 0.000444841f
cc_138 N_GCLKN_14 N_MH_31 0.000153779f
cc_139 N_GCLKN_14 N_MH_33 0.000487925f
cc_140 N_GCLKN_14 N_MM12_g 0.000299262f
cc_141 N_GCLKN_15 N_MM12_g 0.0111767f
cc_142 N_GCLKN_17 N_MH_26 0.000370489f
cc_143 N_GCLKN_5 N_MM12_g 0.000400335f
cc_144 N_GCLKN_3 N_MM0_g 0.000409325f
cc_145 N_GCLKN_20 N_MH_33 0.000475084f
cc_146 N_GCLKN_4 N_MH_27 0.00181763f
cc_147 N_GCLKN_1 N_MH_3 0.00240541f
cc_148 N_GCLKN_17 N_MH_33 0.00132769f
cc_149 N_GCLKN_19 N_MH_33 0.00257615f
cc_150 N_GCLKN_17 N_MH_27 0.00978906f
cc_151 N_MM24_g N_MM12_g 0.0170879f
cc_152 N_GCLKN_14 N_MM0_g 0.0253327f
x_PM_ICGx1_ASAP7_75t_R%CLKN VSS N_MM10_g N_MM20_d N_MM21_d N_CLKN_10 N_CLKN_17
+ N_CLKN_12 N_CLKN_3 N_CLKN_14 N_CLKN_1 N_CLKN_13 N_CLKN_11 N_CLKN_16 N_CLKN_15
+ N_CLKN_4 PM_ICGx1_ASAP7_75t_R%CLKN
cc_153 N_CLKN_10 N_CLK_21 0.000370308f
cc_154 N_CLKN_17 N_CLK_20 0.000263985f
cc_155 N_CLKN_12 N_CLK_15 0.0040314f
cc_156 N_CLKN_3 N_CLK_16 0.000285932f
cc_157 N_CLKN_14 N_CLK_15 0.000297789f
cc_158 N_CLKN_1 N_CLK_8 0.000315502f
cc_159 N_CLKN_13 N_CLK_16 0.00501337f
cc_160 N_CLKN_1 N_CLK_1 0.00141125f
cc_161 N_CLKN_11 N_MM21_g 0.0157643f
cc_162 N_CLKN_16 N_CLK_17 0.000481513f
cc_163 N_CLKN_14 N_CLK_23 0.000517632f
cc_164 N_CLKN_13 N_CLK_23 0.000698225f
cc_165 N_CLKN_15 N_CLK_16 0.00093557f
cc_166 N_CLKN_3 N_MM21_g 0.00094502f
cc_167 N_CLKN_3 N_CLK_3 0.000965282f
cc_168 N_CLKN_4 N_MM21_g 0.00135352f
cc_169 N_CLKN_1 N_CLK_2 0.00148112f
cc_170 N_MM10_g N_MM1_g 0.00161506f
cc_171 N_CLKN_11 N_CLK_3 0.0016435f
cc_172 N_CLKN_16 N_CLK_21 0.00174329f
cc_173 N_MM10_g N_MM9_g 0.00910111f
cc_174 N_CLKN_17 N_CLK_23 0.0259652f
cc_175 N_CLKN_10 N_MM21_g 0.0541698f
x_PM_ICGx1_ASAP7_75t_R%CLK VSS CLK N_MM1_g N_MM9_g N_MM21_g N_MM16_g N_MM13_g
+ N_CLK_23 N_CLK_1 N_CLK_15 N_CLK_21 N_CLK_20 N_CLK_16 N_CLK_8 N_CLK_17 N_CLK_3
+ N_CLK_2 N_CLK_19 N_CLK_22 N_CLK_4 N_CLK_18 PM_ICGx1_ASAP7_75t_R%CLK
cc_176 N_CLK_23 N_NET0121_14 0.0006481f
cc_177 N_CLK_1 N_NET0121_1 0.00164214f
cc_178 N_MM1_g N_MM3_g 0.00327226f
cc_179 N_CLK_15 N_NET0121_14 0.0045553f
x_PM_ICGx1_ASAP7_75t_R%MH VSS N_MM7_g N_MM0_g N_MM12_g N_MM4_d N_MM9_d N_MM1_d
+ N_MM10_d N_MH_23 N_MH_21 N_MH_7 N_MH_19 N_MH_29 N_MH_17 N_MH_27 N_MH_32
+ N_MH_33 N_MH_18 N_MH_3 N_MH_1 N_MH_25 N_MH_26 N_MH_20 N_MH_22 N_MH_24 N_MH_16
+ N_MH_8 N_MH_2 N_MH_30 N_MH_31 PM_ICGx1_ASAP7_75t_R%MH
cc_180 N_MH_23 N_CLK_19 7.89975e-20
cc_181 N_MH_21 N_MM9_g 0.000124493f
cc_182 N_MH_7 N_CLK_15 0.00084646f
cc_183 N_MH_19 N_MM1_g 0.00014953f
cc_184 N_MH_29 N_CLK_19 0.000152172f
cc_185 N_MH_17 N_MM9_g 0.000175721f
cc_186 N_MH_27 N_CLK_22 0.000201848f
cc_187 N_MH_7 N_CLK_1 0.000217949f
cc_188 N_MH_32 N_CLK_16 0.00306034f
cc_189 N_MH_33 N_CLK_4 0.00025201f
cc_190 N_MH_18 N_MM1_g 0.0338858f
cc_191 N_MH_3 N_CLK_4 0.000266711f
cc_192 N_MH_1 N_CLK_8 0.000271258f
cc_193 N_MH_1 N_CLK_20 0.000305803f
cc_194 N_MH_25 N_CLK_20 0.00476157f
cc_195 N_MH_26 N_CLK_16 0.00036254f
cc_196 N_MH_27 N_CLK_4 0.000401496f
cc_197 N_MH_20 N_CLK_15 0.000489331f
cc_198 N_MH_22 N_CLK_8 0.00250131f
cc_199 N_MM7_g N_CLK_8 0.00054433f
cc_200 N_MH_18 N_CLK_1 0.000571045f
cc_201 N_MH_3 N_MM13_g 0.00059973f
cc_202 N_MH_24 N_CLK_23 0.000709745f
cc_203 N_MH_16 N_CLK_2 0.000888436f
cc_204 N_MH_8 N_MM9_g 0.000996974f
cc_205 N_MH_7 N_MM1_g 0.00117547f
cc_206 N_MH_2 N_CLK_3 0.00305765f
cc_207 N_MH_25 N_CLK_19 0.00140162f
cc_208 N_MH_32 N_CLK_17 0.00148652f
cc_209 N_MM12_g N_CLK_4 0.00166619f
cc_210 N_MM0_g N_MM21_g 0.00166641f
cc_211 N_MH_25 N_CLK_23 0.00227901f
cc_212 N_MH_27 N_CLK_18 0.00377115f
cc_213 N_MH_22 N_CLK_19 0.00389174f
cc_214 N_MM12_g N_MM13_g 0.00717608f
cc_215 N_MM0_g N_MM16_g 0.00886723f
cc_216 N_MH_16 N_MM9_g 0.0366524f
cc_217 N_MM0_g N_MM10_g 0.000126632f
cc_218 N_MH_27 N_MM10_g 7.4147e-20
cc_219 N_MM7_g N_MM10_g 9.38753e-20
cc_220 N_MH_17 N_MM10_g 0.000144983f
cc_221 N_MH_32 N_CLKN_15 0.000149897f
cc_222 N_MH_8 N_CLKN_12 0.000161319f
cc_223 N_MH_19 N_MM10_g 0.000166264f
cc_224 N_MH_7 N_CLKN_14 0.000193659f
cc_225 N_MH_30 N_CLKN_14 0.000197641f
cc_226 N_MH_26 N_CLKN_15 0.000214979f
cc_227 N_MH_25 N_CLKN_13 0.000249005f
cc_228 N_MH_24 N_CLKN_3 0.00111962f
cc_229 N_MH_18 N_MM10_g 0.0166804f
cc_230 N_MH_21 N_CLKN_12 0.000497231f
cc_231 N_MH_20 N_CLKN_14 0.00477637f
cc_232 N_MH_23 N_CLKN_14 0.000541328f
cc_233 N_MH_8 N_CLKN_1 0.000680012f
cc_234 N_MH_29 N_CLKN_14 0.000808856f
cc_235 N_MH_8 N_MM10_g 0.00128518f
cc_236 N_MH_7 N_MM10_g 0.0014216f
cc_237 N_MH_16 N_CLKN_1 0.00148339f
cc_238 N_MH_25 N_CLKN_17 0.00330124f
cc_239 N_MH_24 N_CLKN_15 0.00436118f
cc_240 N_MH_22 N_CLKN_12 0.00479639f
cc_241 N_MH_16 N_MM10_g 0.0536123f
cc_242 N_MH_8 N_MM11_g 0.000205147f
cc_243 N_MH_24 N_MM11_g 0.000315363f
cc_244 N_MH_1 N_MS_4 0.00197807f
cc_245 N_MM7_g N_MS_1 0.000552093f
cc_246 N_MH_24 N_MS_1 0.000727436f
cc_247 N_MH_1 N_MS_11 0.0012631f
cc_248 N_MH_22 N_MS_12 0.00131841f
cc_249 N_MH_25 N_MS_13 0.00138738f
cc_250 N_MM7_g N_MS_3 0.00170061f
cc_251 N_MH_25 N_MS_14 0.00239907f
cc_252 N_MM7_g N_MS_10 0.00643105f
cc_253 N_MM7_g N_MS_11 0.00675895f
cc_254 N_MH_24 N_MS_12 0.00369096f
cc_255 N_MH_24 N_MS_15 0.00539925f
cc_256 N_MM7_g N_MM11_g 0.0297006f
*END of ICGx1_ASAP7_75t_R.pxi
.ENDS
** Design:	ICGx2_ASAP7_75t_R
* Created:	"Fri Aug 17 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "ICGx2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "ICGx2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_ICGx2_ASAP7_75t_R%NOS1 VSS 2 3 1
c1 1 VSS 0.000878845f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2160 $X2=0.1080 $Y2=0.2160
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2160 $X2=0.1080 $Y2=0.2160
.ends

.subckt PM_ICGx2_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.0320385f
.ends

.subckt PM_ICGx2_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.00478643f
.ends

.subckt PM_ICGx2_ASAP7_75t_R%SE VSS 8 3 1 4
c1 1 VSS 0.00628739f
c2 3 VSS 0.0830151f
c3 4 VSS 0.00450198f
r1 9 10 2.3902 $w=1.3e-08 $l=1.03e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1267 $X2=0.1350 $Y2=0.1370
r2 8 9 0.408082 $w=1.3e-08 $l=1.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1250 $X2=0.1350 $Y2=0.1267
r3 8 4 6.47102 $w=1.3e-08 $l=2.78e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1250 $X2=0.1350 $Y2=0.0972
r4 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r5 1 10 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1370
.ends

.subckt PM_ICGx2_ASAP7_75t_R%ENA VSS 8 3 1 4
c1 1 VSS 0.00211069f
c2 3 VSS 0.0329546f
c3 4 VSS 0.0100094f
r1 9 10 2.3902 $w=1.3e-08 $l=1.03e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1267 $X2=0.0810 $Y2=0.1370
r2 8 9 0.408082 $w=1.3e-08 $l=1.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1250 $X2=0.0810 $Y2=0.1267
r3 8 4 6.47102 $w=1.3e-08 $l=2.78e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1250 $X2=0.0810 $Y2=0.0972
r4 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r5 1 10 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1370
.ends

.subckt PM_ICGx2_ASAP7_75t_R%noxref_26 VSS 1
c1 1 VSS 0.0423594f
.ends

.subckt PM_ICGx2_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.0423312f
.ends

.subckt PM_ICGx2_ASAP7_75t_R%GCLK VSS 22 16 17 30 31 7 8 11 1 2 10 9
c1 1 VSS 0.0100082f
c2 2 VSS 0.0101158f
c3 7 VSS 0.00460999f
c4 8 VSS 0.00453219f
c5 9 VSS 0.011605f
c6 10 VSS 0.00918593f
c7 11 VSS 0.00744682f
c8 12 VSS 0.00335907f
c9 13 VSS 0.00352401f
r1 31 29 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9350 $Y=0.2025 $X2=0.9325 $Y2=0.2025
r2 2 29 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9180 $Y=0.2025 $X2=0.9325 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9035 $Y=0.2025 $X2=0.9180 $Y2=0.2025
r4 30 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9010 $Y=0.2025 $X2=0.9035 $Y2=0.2025
r5 2 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.9180 $Y=0.2025
+ $X2=0.9180 $Y2=0.2340
r6 25 26 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.2340 $X2=0.9585 $Y2=0.2340
r7 10 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.9045
+ $Y=0.2340 $X2=0.9180 $Y2=0.2340
r8 13 24 2.6649 $w=1.77676e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9990 $Y=0.2340 $X2=0.9990 $Y2=0.2155
r9 13 26 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9990 $Y=0.2340 $X2=0.9585 $Y2=0.2340
r10 23 24 6.8208 $w=1.3e-08 $l=2.93e-08 $layer=M1 $thickness=3.6e-08 $X=0.9990
+ $Y=0.1862 $X2=0.9990 $Y2=0.2155
r11 22 23 4.72209 $w=1.3e-08 $l=2.02e-08 $layer=M1 $thickness=3.6e-08 $X=0.9990
+ $Y=0.1660 $X2=0.9990 $Y2=0.1862
r12 22 21 12.0676 $w=1.3e-08 $l=5.18e-08 $layer=M1 $thickness=3.6e-08 $X=0.9990
+ $Y=0.1660 $X2=0.9990 $Y2=0.1142
r13 11 12 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.9990
+ $Y=0.0540 $X2=0.9990 $Y2=0.0360
r14 11 21 14.0497 $w=1.3e-08 $l=6.02e-08 $layer=M1 $thickness=3.6e-08 $X=0.9990
+ $Y=0.0540 $X2=0.9990 $Y2=0.1142
r15 12 20 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9990 $Y=0.0360 $X2=0.9585 $Y2=0.0360
r16 19 20 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.0360 $X2=0.9585 $Y2=0.0360
r17 18 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.9045
+ $Y=0.0360 $X2=0.9180 $Y2=0.0360
r18 9 18 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.8895
+ $Y=0.0360 $X2=0.9045 $Y2=0.0360
r19 1 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.9180 $Y=0.0675
+ $X2=0.9180 $Y2=0.0360
r20 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9350 $Y=0.0675 $X2=0.9325 $Y2=0.0675
r21 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9180 $Y=0.0675 $X2=0.9325 $Y2=0.0675
r22 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9035 $Y=0.0675 $X2=0.9180 $Y2=0.0675
r23 16 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9010 $Y=0.0675 $X2=0.9035 $Y2=0.0675
.ends

.subckt PM_ICGx2_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.00366067f
.ends

.subckt PM_ICGx2_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.00364721f
.ends

.subckt PM_ICGx2_ASAP7_75t_R%NET0121 VSS 9 41 42 44 11 13 4 3 12 10 1 14
c1 1 VSS 0.00374778f
c2 3 VSS 0.0071602f
c3 4 VSS 0.0090272f
c4 9 VSS 0.0801723f
c5 10 VSS 0.00629634f
c6 11 VSS 0.00495902f
c7 12 VSS 0.0168136f
c8 13 VSS 0.0104772f
c9 14 VSS 0.0067057f
c10 15 VSS 0.00312965f
c11 16 VSS 0.00353835f
r1 44 43 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r2 11 43 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r3 42 40 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0540 $X2=0.1225 $Y2=0.0540
r4 4 40 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0540 $X2=0.1225 $Y2=0.0540
r5 10 4 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0540 $X2=0.1080 $Y2=0.0540
r6 41 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0540 $X2=0.0935 $Y2=0.0540
r7 3 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0540 $Y2=0.2330
r8 4 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0540
+ $X2=0.1080 $Y2=0.0360
r9 37 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2330 $X2=0.0675 $Y2=0.2330
r10 35 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.2330 $X2=0.0675 $Y2=0.2330
r11 34 35 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2330 $X2=0.0810 $Y2=0.2330
r12 33 34 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2330 $X2=0.1080 $Y2=0.2330
r13 12 16 5.06479 $w=1.46038e-08 $l=2.70046e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1620 $Y=0.2330 $X2=0.1890 $Y2=0.2325
r14 12 33 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2330 $X2=0.1350 $Y2=0.2330
r15 30 31 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.1215 $Y2=0.0360
r16 28 31 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1215 $Y2=0.0360
r17 13 15 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1620 $Y=0.0360 $X2=0.1890 $Y2=0.0360
r18 13 28 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r19 16 26 0.983973 $w=1.77222e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2325 $X2=0.1890 $Y2=0.2235
r20 15 21 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1890 $Y2=0.0575
r21 25 26 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2110 $X2=0.1890 $Y2=0.2235
r22 24 25 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1985 $X2=0.1890 $Y2=0.2110
r23 23 24 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1910 $X2=0.1890 $Y2=0.1985
r24 22 23 9.211 $w=1.3e-08 $l=3.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1515 $X2=0.1890 $Y2=0.1910
r25 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0710 $X2=0.1890 $Y2=0.0575
r26 19 20 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0810 $X2=0.1890 $Y2=0.0710
r27 14 19 5.47996 $w=1.3e-08 $l=2.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1045 $X2=0.1890 $Y2=0.0810
r28 14 22 10.9599 $w=1.3e-08 $l=4.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1045 $X2=0.1890 $Y2=0.1515
r29 9 1 6.2219 $w=1.2115e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1340
r30 1 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1340
+ $X2=0.1890 $Y2=0.1515
r31 3 11 1e-05
.ends

.subckt PM_ICGx2_ASAP7_75t_R%PU1 VSS 5 8 3 1
c1 1 VSS 0.00536697f
c2 3 VSS 0.00340041f
r1 8 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r2 6 7 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2260 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r3 1 6 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2140 $Y=0.2025 $X2=0.2260 $Y2=0.2025
r4 3 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2140 $Y2=0.2025
r5 5 3 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
.ends

.subckt PM_ICGx2_ASAP7_75t_R%PD3 VSS 5 8 3 1
c1 1 VSS 0.00335173f
c2 3 VSS 0.00246874f
r1 8 7 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0405 $X2=0.3925 $Y2=0.0405
r2 1 7 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3800 $Y=0.0405 $X2=0.3925 $Y2=0.0405
r3 4 1 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3680 $Y=0.0405 $X2=0.3800 $Y2=0.0405
r4 3 4 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.0405 $X2=0.3680 $Y2=0.0405
r5 5 3 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0405 $X2=0.3635 $Y2=0.0405
.ends

.subckt PM_ICGx2_ASAP7_75t_R%NET0140 VSS 2 3 1
c1 1 VSS 0.000934541f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.0675 $X2=0.8100 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8270 $Y=0.0675 $X2=0.8100 $Y2=0.0675
.ends

.subckt PM_ICGx2_ASAP7_75t_R%PD1 VSS 7 10 4 5 1
c1 1 VSS 0.0097948f
c2 4 VSS 0.00323902f
c3 5 VSS 0.00185993f
r1 10 9 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r2 8 9 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2800 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r3 5 8 0.123457 $w=8.1e-08 $l=1e-08 $layer=N_src_drn $thickness=1e-09 $X=0.2700
+ $Y=0.0675 $X2=0.2800 $Y2=0.0675
r4 4 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0675 $X2=0.2140 $Y2=0.0675
r5 7 4 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2015 $Y2=0.0675
r6 1 5 1e-05
.ends

.subckt PM_ICGx2_ASAP7_75t_R%NET0141 VSS 2 3 1
c1 1 VSS 0.000863663f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.0675 $X2=0.7020 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.0675 $X2=0.7020 $Y2=0.0675
.ends

.subckt PM_ICGx2_ASAP7_75t_R%PD2 VSS 7 13 5 4 1
c1 1 VSS 0.00729312f
c2 4 VSS 0.00188002f
c3 5 VSS 0.0023855f
r1 13 12 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r2 5 12 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3800 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r3 10 5 9.87715 $w=2.32e-08 $l=2.1e-08 $layer=LISD $thickness=2.7e-08 $X=0.3570
+ $Y=0.2295 $X2=0.3780 $Y2=0.2295
r4 9 10 6.11443 $w=2.32e-08 $l=1.3e-08 $layer=LISD $thickness=2.7e-08 $X=0.3440
+ $Y=0.2295 $X2=0.3570 $Y2=0.2295
r5 8 9 2.82204 $w=2.32e-08 $l=6e-09 $layer=LISD $thickness=2.7e-08 $X=0.3380
+ $Y=0.2295 $X2=0.3440 $Y2=0.2295
r6 1 8 6.58477 $w=2.32e-08 $l=1.4e-08 $layer=LISD $thickness=2.7e-08 $X=0.3240
+ $Y=0.2295 $X2=0.3380 $Y2=0.2295
r7 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2295 $X2=0.3220 $Y2=0.2295
r8 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2295 $X2=0.3095 $Y2=0.2295
.ends

.subckt PM_ICGx2_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.00441216f
.ends

.subckt PM_ICGx2_ASAP7_75t_R%GCLKN VSS 12 13 50 51 59 60 63 64 14 5 15 3 17 4
+ 16 18 21 1 20 23 22
c1 1 VSS 0.00744186f
c2 3 VSS 0.0084736f
c3 4 VSS 0.00526014f
c4 5 VSS 0.00812327f
c5 12 VSS 0.0806139f
c6 13 VSS 0.0809716f
c7 14 VSS 0.00482359f
c8 15 VSS 0.00542911f
c9 16 VSS 0.00541249f
c10 17 VSS 0.0130726f
c11 18 VSS 0.00673268f
c12 19 VSS 0.0016096f
c13 20 VSS 0.00288977f
c14 21 VSS 0.00387804f
c15 22 VSS 0.000552432f
c16 23 VSS 0.000847186f
r1 64 62 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.2160 $X2=0.7165 $Y2=0.2160
r2 3 62 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7020 $Y=0.2160 $X2=0.7165 $Y2=0.2160
r3 15 3 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.2160 $X2=0.7020 $Y2=0.2160
r4 63 15 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.2160 $X2=0.6875 $Y2=0.2160
r5 60 58 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8270 $Y=0.2160 $X2=0.8245 $Y2=0.2160
r6 5 58 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8100 $Y=0.2160 $X2=0.8245 $Y2=0.2160
r7 16 5 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.2160 $X2=0.8100 $Y2=0.2160
r8 59 16 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.2160 $X2=0.7955 $Y2=0.2160
r9 3 55 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7020 $Y=0.2160
+ $X2=0.7020 $Y2=0.2310
r10 5 52 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8100 $Y=0.2160
+ $X2=0.8100 $Y2=0.2310
r11 55 56 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.2310 $X2=0.7380 $Y2=0.2310
r12 52 53 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.2310 $X2=0.8235 $Y2=0.2310
r13 17 52 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.2310 $X2=0.8100 $Y2=0.2310
r14 17 56 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.2310 $X2=0.7380 $Y2=0.2310
r15 50 49 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.0675 $X2=0.7705 $Y2=0.0675
r16 4 49 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7560 $Y=0.0675 $X2=0.7705 $Y2=0.0675
r17 14 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7415 $Y=0.0675 $X2=0.7560 $Y2=0.0675
r18 51 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.0675 $X2=0.7415 $Y2=0.0675
r19 46 53 1.20242 $w=1.425e-08 $l=1.54434e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8370 $Y=0.2235 $X2=0.8235 $Y2=0.2310
r20 45 46 2.01858 $w=1.37895e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.8370 $Y=0.2140 $X2=0.8370 $Y2=0.2235
r21 44 45 2.37574 $w=1.49231e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8370 $Y=0.2010 $X2=0.8370 $Y2=0.2140
r22 21 44 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1920 $X2=0.8370 $Y2=0.2010
r23 4 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7560 $Y=0.0675
+ $X2=0.7560 $Y2=0.0720
r24 19 23 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8640 $Y=0.1970 $X2=0.8910 $Y2=0.1970
r25 19 21 4.60559 $w=1.39091e-08 $l=2.74591e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8640 $Y=0.1970 $X2=0.8370 $Y2=0.1920
r26 42 43 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.0720 $X2=0.7965 $Y2=0.0720
r27 40 43 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.0720 $X2=0.7965 $Y2=0.0720
r28 39 40 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.8625
+ $Y=0.0720 $X2=0.8370 $Y2=0.0720
r29 18 22 0.79938 $w=1.72857e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8805 $Y=0.0720 $X2=0.8910 $Y2=0.0720
r30 18 39 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8805
+ $Y=0.0720 $X2=0.8625 $Y2=0.0720
r31 23 37 5.22999 $w=1.59898e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8910 $Y=0.1970 $X2=0.8910 $Y2=0.1675
r32 22 36 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.0720 $X2=0.8910 $Y2=0.0900
r33 13 32 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=0.9450
+ $Y=0.1350 $X2=0.9450 $Y2=0.1360
r34 35 37 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1460 $X2=0.8910 $Y2=0.1675
r35 34 35 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1360 $X2=0.8910 $Y2=0.1460
r36 20 34 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1130 $X2=0.8910 $Y2=0.1360
r37 20 36 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1130 $X2=0.8910 $Y2=0.0900
r38 30 32 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9325 $Y=0.1360 $X2=0.9450 $Y2=0.1360
r39 29 30 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9180 $Y=0.1360 $X2=0.9325 $Y2=0.1360
r40 28 29 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9035 $Y=0.1360 $X2=0.9180 $Y2=0.1360
r41 26 28 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.9005 $Y=0.1360 $X2=0.9035 $Y2=0.1360
r42 25 26 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.8910
+ $Y=0.1360 $X2=0.9005 $Y2=0.1360
r43 25 34 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8910 $Y=0.1360
+ $X2=0.8910 $Y2=0.1360
r44 1 25 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.8815
+ $Y=0.1360 $X2=0.8910 $Y2=0.1360
r45 1 27 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.8815
+ $Y=0.1360 $X2=0.8805 $Y2=0.1360
r46 12 25 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.8910 $Y=0.1350 $X2=0.8910 $Y2=0.1360
r47 12 27 0.610027 $w=2.16919e-07 $l=1.05475e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.8910 $Y=0.1350 $X2=0.8805 $Y2=0.1360
r48 12 28 1.79147 $w=1.8466e-07 $l=1.25399e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.8910 $Y=0.1350 $X2=0.9035 $Y2=0.1360
.ends

.subckt PM_ICGx2_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.00423341f
.ends

.subckt PM_ICGx2_ASAP7_75t_R%CLK VSS 49 10 11 12 13 14 23 1 15 21 20 16 8 17 3
+ 2 19 22 4 18
c1 1 VSS 0.0038099f
c2 2 VSS 0.00185515f
c3 3 VSS 0.00735746f
c4 4 VSS 0.00894294f
c5 8 VSS 0.00398121f
c6 10 VSS 0.00630487f
c7 11 VSS 0.00625709f
c8 12 VSS 0.0820738f
c9 13 VSS 0.034238f
c10 14 VSS 0.0342767f
c11 15 VSS 0.00470944f
c12 16 VSS 0.00460581f
c13 17 VSS 0.00487152f
c14 18 VSS 0.0022609f
c15 19 VSS 0.00194584f
c16 20 VSS 0.00384565f
c17 21 VSS 0.00245608f
c18 22 VSS 0.00241574f
c19 23 VSS 0.00589905f
r1 2 78 3.16825 $w=2.1e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.3520
+ $Y=0.1335 $X2=0.3555 $Y2=0.1335
r2 11 2 3.48292 $w=1.19095e-07 $l=1.80278e-09 $layer=LIG $thickness=5.18095e-08
+ $X=0.3510 $Y=0.1350 $X2=0.3520 $Y2=0.1335
r3 77 78 4.91375 $w=2.12e-08 $l=1.5e-09 $layer=LISD $thickness=2.7e-08
+ $X=0.3570 $Y=0.1335 $X2=0.3555 $Y2=0.1335
r4 76 77 11.4654 $w=2.12e-08 $l=2.1e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.3780 $Y=0.1335 $X2=0.3570 $Y2=0.1335
r5 75 76 7.37062 $w=2.12e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.3915 $Y=0.1335 $X2=0.3780 $Y2=0.1335
r6 8 73 5.7327 $w=2.12e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08 $X=0.3945
+ $Y=0.1335 $X2=0.4050 $Y2=0.1335
r7 8 75 1.63792 $w=2.12e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.3945
+ $Y=0.1335 $X2=0.3915 $Y2=0.1335
r8 1 62 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1335
+ $X2=0.2430 $Y2=0.1330
r9 10 1 3.19489 $w=1.24e-07 $l=1.5e-09 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1335
r10 69 70 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1340 $X2=0.4050 $Y2=0.1435
r11 69 73 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4050 $Y=0.1340
+ $X2=0.4050 $Y2=0.1335
r12 19 20 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1530 $X2=0.4230 $Y2=0.1530
r13 19 70 1.03499 $w=1.77368e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.1530 $X2=0.4050 $Y2=0.1435
r14 63 64 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1430 $X2=0.2430 $Y2=0.1530
r15 62 63 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1330 $X2=0.2430 $Y2=0.1430
r16 15 62 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1215 $X2=0.2430 $Y2=0.1330
r17 20 54 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4230 $Y=0.1530
+ $X2=0.4230 $Y2=0.1530
r18 3 46 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6210 $Y=0.1350
+ $X2=0.6210 $Y2=0.1330
r19 12 3 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1350
r20 57 58 7.22888 $w=1.3e-08 $l=3.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1530 $X2=0.2740 $Y2=0.1530
r21 57 64 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.2430 $Y=0.1530
+ $X2=0.2430 $Y2=0.1530
r22 54 55 19.5879 $w=1.3e-08 $l=8.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.4230
+ $Y=0.1530 $X2=0.5070 $Y2=0.1530
r23 53 54 15.8569 $w=1.3e-08 $l=6.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.3550
+ $Y=0.1530 $X2=0.4230 $Y2=0.1530
r24 53 58 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.3550
+ $Y=0.1530 $X2=0.2740 $Y2=0.1530
r25 50 51 5.07188 $w=1.3e-08 $l=2.18e-08 $layer=M2 $thickness=3.6e-08 $X=0.5992
+ $Y=0.1530 $X2=0.6210 $Y2=0.1530
r26 49 50 3.08976 $w=1.3e-08 $l=1.32e-08 $layer=M2 $thickness=3.6e-08 $X=0.5860
+ $Y=0.1530 $X2=0.5992 $Y2=0.1530
r27 49 23 0.524677 $w=1.3e-08 $l=2.3e-09 $layer=M2 $thickness=3.6e-08 $X=0.5860
+ $Y=0.1530 $X2=0.5837 $Y2=0.1530
r28 23 55 17.8973 $w=1.3e-08 $l=7.67e-08 $layer=M2 $thickness=3.6e-08 $X=0.5837
+ $Y=0.1530 $X2=0.5070 $Y2=0.1530
r29 47 48 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1430 $X2=0.6210 $Y2=0.1455
r30 46 47 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1330 $X2=0.6210 $Y2=0.1430
r31 16 44 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1545 $X2=0.6210 $Y2=0.1700
r32 16 48 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1545 $X2=0.6210 $Y2=0.1455
r33 16 51 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.6210 $Y=0.1545
+ $X2=0.6210 $Y2=0.1530
r34 21 43 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.1870 $X2=0.6480 $Y2=0.1870
r35 21 44 2.31511 $w=1.81882e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.1870 $X2=0.6210 $Y2=0.1700
r36 42 43 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1870 $X2=0.6480 $Y2=0.1870
r37 41 42 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6860
+ $Y=0.1870 $X2=0.6750 $Y2=0.1870
r38 17 22 7.38932 $w=1.37246e-08 $l=3.87072e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7175 $Y=0.1870 $X2=0.7560 $Y2=0.1830
r39 17 41 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.7175
+ $Y=0.1870 $X2=0.6860 $Y2=0.1870
r40 22 38 1.32639 $w=1.59412e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.7560 $Y=0.1830 $X2=0.7560 $Y2=0.1745
r41 13 33 2.92627 $w=1.245e-07 $l=2.7e-08 $layer=LIG $thickness=5.2e-08
+ $X=0.7290 $Y=0.1350 $X2=0.7290 $Y2=0.1620
r42 37 38 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.1620 $X2=0.7560 $Y2=0.1745
r43 36 37 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.1500 $X2=0.7560 $Y2=0.1620
r44 18 36 1.28254 $w=1.3e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.1445 $X2=0.7560 $Y2=0.1500
r45 31 33 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7415 $Y=0.1620 $X2=0.7290 $Y2=0.1620
r46 30 31 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7560 $Y=0.1620 $X2=0.7415 $Y2=0.1620
r47 30 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7560 $Y=0.1620
+ $X2=0.7560 $Y2=0.1620
r48 29 30 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7705 $Y=0.1620 $X2=0.7560 $Y2=0.1620
r49 4 28 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.7830
+ $Y=0.1620 $X2=0.7830 $Y2=0.1620
r50 4 29 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7830 $Y=0.1620 $X2=0.7705 $Y2=0.1620
r51 4 35 2.90696 $w=2.1681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7830 $Y=0.1620 $X2=0.7935 $Y2=0.1620
r52 28 29 1.47681 $w=1.53e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7830 $Y=0.1620 $X2=0.7705 $Y2=0.1620
r53 28 35 0.295362 $w=1.53e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7830 $Y=0.1620 $X2=0.7935 $Y2=0.1620
r54 14 28 0.314665 $w=2.27e-07 $l=2.7e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.7830 $Y=0.1350 $X2=0.7830 $Y2=0.1620
.ends

.subckt PM_ICGx2_ASAP7_75t_R%MS VSS 9 40 46 1 12 13 15 3 14 4 11 10
c1 1 VSS 0.00207793f
c2 3 VSS 0.0050376f
c3 4 VSS 0.00604156f
c4 9 VSS 0.0369211f
c5 10 VSS 0.00306725f
c6 11 VSS 0.00310605f
c7 12 VSS 0.00122497f
c8 13 VSS 0.00124628f
c9 14 VSS 0.00665953f
c10 15 VSS 0.000349834f
r1 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2295 $X2=0.4840 $Y2=0.2295
r2 46 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2295 $X2=0.4715 $Y2=0.2295
r3 4 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2295
+ $X2=0.4860 $Y2=0.2330
r4 42 43 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.2330 $X2=0.4990 $Y2=0.2330
r5 14 38 1.06916 $w=1.78e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.2330 $X2=0.5125 $Y2=0.2235
r6 14 43 1.90218 $w=1.65185e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5125 $Y=0.2330 $X2=0.4990 $Y2=0.2330
r7 10 31 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0405 $X2=0.4840 $Y2=0.0405
r8 40 10 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0405 $X2=0.4715 $Y2=0.0405
r9 37 38 2.49333 $w=1.4e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.2110 $X2=0.5125 $Y2=0.2235
r10 36 37 4.1888 $w=1.4e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.1900 $X2=0.5125 $Y2=0.2110
r11 35 36 3.69013 $w=1.4e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.1715 $X2=0.5125 $Y2=0.1900
r12 34 35 3.69013 $w=1.4e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.1530 $X2=0.5125 $Y2=0.1715
r13 33 34 4.1888 $w=1.4e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.1320 $X2=0.5125 $Y2=0.1530
r14 32 33 4.88693 $w=1.4e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.1075 $X2=0.5125 $Y2=0.1320
r15 13 15 0.843012 $w=1.80909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5125 $Y=0.0930 $X2=0.5125 $Y2=0.0820
r16 13 32 2.89227 $w=1.4e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.0930 $X2=0.5125 $Y2=0.1075
r17 3 29 10.904 $w=2.02e-08 $l=1.85e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4860 $Y=0.0635 $X2=0.4860 $Y2=0.0820
r18 3 31 13.5563 $w=2.02e-08 $l=2.3e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4860 $Y=0.0635 $X2=0.4860 $Y2=0.0405
r19 15 28 1.37684 $w=2.03185e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5125 $Y=0.0820 $X2=0.4990 $Y2=0.0820
r20 27 28 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.0820 $X2=0.4990 $Y2=0.0820
r21 27 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0820
+ $X2=0.4860 $Y2=0.0820
r22 26 27 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4750
+ $Y=0.0820 $X2=0.4860 $Y2=0.0820
r23 25 26 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4600
+ $Y=0.0820 $X2=0.4750 $Y2=0.0820
r24 24 25 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4310
+ $Y=0.0820 $X2=0.4600 $Y2=0.0820
r25 23 24 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.4145
+ $Y=0.0820 $X2=0.4310 $Y2=0.0820
r26 21 23 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4055
+ $Y=0.0820 $X2=0.4145 $Y2=0.0820
r27 12 21 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3965
+ $Y=0.0820 $X2=0.4055 $Y2=0.0820
r28 18 20 2.94116 $w=2.133e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.4060
+ $Y=0.0820 $X2=0.4160 $Y2=0.0820
r29 18 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4060 $Y=0.0820
+ $X2=0.4055 $Y2=0.0820
r30 1 18 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.3960
+ $Y=0.0820 $X2=0.4060 $Y2=0.0820
r31 1 19 0.851883 $w=1.865e-08 $l=2e-09 $layer=LIG $thickness=4.8e-08 $X=0.3960
+ $Y=0.0820 $X2=0.3940 $Y2=0.0820
r32 17 18 2.35044 $w=2.2e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.4050
+ $Y=0.0820 $X2=0.4060 $Y2=0.0820
r33 17 19 0.590723 $w=1.53e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4050 $Y=0.0820 $X2=0.3940 $Y2=0.0820
r34 17 20 0.590723 $w=1.53e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4050 $Y=0.0820 $X2=0.4160 $Y2=0.0820
r35 9 17 0.314665 $w=2.27e-07 $l=5.3e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4050 $Y2=0.0820
.ends

.subckt PM_ICGx2_ASAP7_75t_R%CLKN VSS 9 53 55 10 13 18 3 15 12 1 17 11 14 16 4
c1 1 VSS 0.000101024f
c2 3 VSS 0.00618941f
c3 4 VSS 0.00785619f
c4 9 VSS 0.00447201f
c5 10 VSS 0.00630299f
c6 11 VSS 0.00632934f
c7 12 VSS 0.000537869f
c8 13 VSS 0.00123396f
c9 14 VSS 0.00264632f
c10 15 VSS 0.000650934f
c11 16 VSS 0.000859628f
c12 17 VSS 0.00632012f
c13 18 VSS 0.00922488f
r1 55 54 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.2025 $X2=0.6085 $Y2=0.2025
r2 11 54 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5960 $Y=0.2025 $X2=0.6085 $Y2=0.2025
r3 53 52 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.0675 $X2=0.6085 $Y2=0.0675
r4 10 52 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5960 $Y=0.0675 $X2=0.6085 $Y2=0.0675
r5 4 46 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2295
+ $X2=0.5940 $Y2=0.2320
r6 3 43 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0605
+ $X2=0.5940 $Y2=0.0860
r7 45 46 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5810
+ $Y=0.2320 $X2=0.5940 $Y2=0.2320
r8 17 41 1.03499 $w=1.77368e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.5680 $Y=0.2320 $X2=0.5680 $Y2=0.2225
r9 17 45 1.85116 $w=1.64615e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5680 $Y=0.2320 $X2=0.5810 $Y2=0.2320
r10 42 43 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5810
+ $Y=0.0860 $X2=0.5940 $Y2=0.0860
r11 16 38 3.36689 $w=1.53077e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5680 $Y=0.0860 $X2=0.5680 $Y2=0.1055
r12 16 42 1.85116 $w=1.64615e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5680 $Y=0.0860 $X2=0.5810 $Y2=0.0860
r13 40 41 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5680
+ $Y=0.2100 $X2=0.5680 $Y2=0.2225
r14 39 40 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5680
+ $Y=0.1970 $X2=0.5680 $Y2=0.2100
r15 37 39 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5680
+ $Y=0.1880 $X2=0.5680 $Y2=0.1970
r16 13 37 9.32759 $w=1.3e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.5680
+ $Y=0.1480 $X2=0.5680 $Y2=0.1880
r17 13 38 9.91056 $w=1.3e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5680
+ $Y=0.1480 $X2=0.5680 $Y2=0.1055
r18 35 37 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.5680 $Y=0.1890
+ $X2=0.5680 $Y2=0.1880
r19 34 35 30.0815 $w=1.3e-08 $l=1.29e-07 $layer=M2 $thickness=3.6e-08 $X=0.4390
+ $Y=0.1890 $X2=0.5680 $Y2=0.1890
r20 33 34 30.0815 $w=1.3e-08 $l=1.29e-07 $layer=M2 $thickness=3.6e-08 $X=0.3100
+ $Y=0.1890 $X2=0.4390 $Y2=0.1890
r21 18 33 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.2985
+ $Y=0.1890 $X2=0.3100 $Y2=0.1890
r22 31 33 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.3145 $Y=0.1890
+ $X2=0.3100 $Y2=0.1890
r23 30 31 1.51573 $w=1.3e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3080
+ $Y=0.1890 $X2=0.3145 $Y2=0.1890
r24 29 30 0.721491 $w=1.57778e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.3035 $Y=0.1890 $X2=0.3080 $Y2=0.1890
r25 15 29 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2945
+ $Y=0.1890 $X2=0.3035 $Y2=0.1890
r26 27 29 4.68572 $w=1.35814e-08 $l=2.87446e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1610 $X2=0.3035 $Y2=0.1890
r27 26 27 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1330 $X2=0.2970 $Y2=0.1610
r28 25 26 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1215 $X2=0.2970 $Y2=0.1330
r29 12 25 3.96423 $w=1.3e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1045 $X2=0.2970 $Y2=0.1215
r30 12 14 4.29965 $w=1.49149e-08 $l=2.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1045 $X2=0.2970 $Y2=0.0810
r31 1 22 2.88023 $w=2.1e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.2970
+ $Y=0.1335 $X2=0.2970 $Y2=0.1335
r32 1 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1335
+ $X2=0.2970 $Y2=0.1330
r33 9 22 0.314665 $w=2.27e-07 $l=1.5e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2970 $Y2=0.1335
r34 4 11 1e-05
r35 3 10 1e-05
.ends

.subckt PM_ICGx2_ASAP7_75t_R%MH VSS 13 14 15 77 81 100 104 23 7 21 29 19 17 27
+ 32 33 18 3 1 25 26 20 22 24 16 8 2 30 31
c1 1 VSS 0.0023512f
c2 2 VSS 0.0046007f
c3 3 VSS 0.00401071f
c4 7 VSS 0.00517367f
c5 8 VSS 0.00493236f
c6 13 VSS 0.036861f
c7 14 VSS 0.0818838f
c8 15 VSS 0.0818348f
c9 16 VSS 0.00317832f
c10 17 VSS 0.000556973f
c11 18 VSS 0.00315327f
c12 19 VSS 0.000592325f
c13 20 VSS 0.00828793f
c14 21 VSS 0.00486108f
c15 22 VSS 0.000832664f
c16 23 VSS 0.000426805f
c17 24 VSS 0.0293109f
c18 25 VSS 0.00200931f
c19 26 VSS 0.00222408f
c20 27 VSS 0.00203078f
c21 28 VSS 0.00226764f
c22 29 VSS 7.47383e-20
c23 30 VSS 0.00263428f
c24 31 VSS 0.00334412f
c25 32 VSS 0.000688482f
c26 33 VSS 0.00130174f
r1 104 103 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2295 $X2=0.2845 $Y2=0.2295
r2 102 103 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2800 $Y=0.2295 $X2=0.2845 $Y2=0.2295
r3 18 102 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2680 $Y=0.2295 $X2=0.2800 $Y2=0.2295
r4 19 18 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2295 $X2=0.2680 $Y2=0.2295
r5 98 99 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.1890 $X2=0.2600 $Y2=0.1890
r6 100 98 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.1890 $X2=0.2555 $Y2=0.1890
r7 18 99 0.185185 $w=5.4e-08 $l=1e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.1890 $X2=0.2600 $Y2=0.1890
r8 7 94 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2295
+ $X2=0.2700 $Y2=0.2320
r9 7 18 23.8708 $w=2.02e-08 $l=4.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.2700 $Y=0.2295 $X2=0.2700 $Y2=0.1890
r10 94 95 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2320 $X2=0.2835 $Y2=0.2320
r11 92 95 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3060
+ $Y=0.2320 $X2=0.2835 $Y2=0.2320
r12 20 30 2.96589 $w=1.31923e-08 $l=2.31193e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3365 $Y=0.2320 $X2=0.3580 $Y2=0.2235
r13 20 92 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.3365
+ $Y=0.2320 $X2=0.3060 $Y2=0.2320
r14 1 86 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1900
+ $X2=0.4590 $Y2=0.1900
r15 13 1 3.49039 $w=1.235e-07 $l=5.5e-08 $layer=LIG $thickness=5.2e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4590 $Y2=0.1900
r16 23 75 2.8493 $w=1.32e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.2110 $X2=0.3580 $Y2=0.1985
r17 23 30 2.8493 $w=1.32e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.2110 $X2=0.3580 $Y2=0.2235
r18 85 86 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4485
+ $Y=0.1900 $X2=0.4590 $Y2=0.1900
r19 84 85 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4305
+ $Y=0.1900 $X2=0.4485 $Y2=0.1900
r20 83 84 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1900 $X2=0.4305 $Y2=0.1900
r21 82 83 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3940
+ $Y=0.1900 $X2=0.4050 $Y2=0.1900
r22 25 29 3.78225 $w=1.50238e-08 $l=2.15058e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3795 $Y=0.1900 $X2=0.3580 $Y2=0.1895
r23 25 82 3.38125 $w=1.3e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3795
+ $Y=0.1900 $X2=0.3940 $Y2=0.1900
r24 81 80 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0405 $X2=0.3385 $Y2=0.0405
r25 79 80 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3340 $Y=0.0405 $X2=0.3385 $Y2=0.0405
r26 8 79 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3220 $Y=0.0405 $X2=0.3340 $Y2=0.0405
r27 17 8 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0405 $X2=0.3220 $Y2=0.0405
r28 16 8 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0810 $X2=0.3220 $Y2=0.0810
r29 77 16 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0810 $X2=0.3095 $Y2=0.0810
r30 29 70 0.983973 $w=1.77222e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.3580 $Y=0.1895 $X2=0.3580 $Y2=0.1805
r31 29 75 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.1895 $X2=0.3580 $Y2=0.1985
r32 8 63 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0405
+ $X2=0.3195 $Y2=0.0360
r33 69 70 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.1710 $X2=0.3580 $Y2=0.1805
r34 68 69 6.99569 $w=1.3e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.1410 $X2=0.3580 $Y2=0.1710
r35 67 68 8.27824 $w=1.3e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.1055 $X2=0.3580 $Y2=0.1410
r36 66 67 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.0905 $X2=0.3580 $Y2=0.1055
r37 65 66 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.0815 $X2=0.3580 $Y2=0.0905
r38 64 65 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.0725 $X2=0.3580 $Y2=0.0815
r39 22 28 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.0585 $X2=0.3580 $Y2=0.0360
r40 22 64 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.0585 $X2=0.3580 $Y2=0.0725
r41 21 61 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3285
+ $Y=0.0360 $X2=0.3410 $Y2=0.0360
r42 21 63 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3285
+ $Y=0.0360 $X2=0.3195 $Y2=0.0360
r43 28 60 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3580 $Y=0.0360 $X2=0.3795 $Y2=0.0360
r44 28 61 2.78392 $w=1.56471e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3580 $Y=0.0360 $X2=0.3410 $Y2=0.0360
r45 59 60 18.0722 $w=1.3e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.4570
+ $Y=0.0360 $X2=0.3795 $Y2=0.0360
r46 58 59 19.4713 $w=1.3e-08 $l=8.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5405
+ $Y=0.0360 $X2=0.4570 $Y2=0.0360
r47 57 58 10.1438 $w=1.3e-08 $l=4.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5840
+ $Y=0.0360 $X2=0.5405 $Y2=0.0360
r48 56 57 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.6105
+ $Y=0.0360 $X2=0.5840 $Y2=0.0360
r49 55 56 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0360 $X2=0.6105 $Y2=0.0360
r50 24 31 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6480 $Y=0.0360 $X2=0.6750 $Y2=0.0360
r51 24 55 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.6480
+ $Y=0.0360 $X2=0.6210 $Y2=0.0360
r52 31 51 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0360 $X2=0.6750 $Y2=0.0540
r53 2 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6750 $Y=0.1350
+ $X2=0.6750 $Y2=0.1330
r54 14 2 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6750
+ $Y=0.1350 $X2=0.6750 $Y2=0.1350
r55 50 51 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0680 $X2=0.6750 $Y2=0.0540
r56 49 50 1.63233 $w=1.3e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0750 $X2=0.6750 $Y2=0.0680
r57 48 49 0.932759 $w=1.3e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0790 $X2=0.6750 $Y2=0.0750
r58 47 48 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0880 $X2=0.6750 $Y2=0.0790
r59 26 32 1.33376 $w=1.70476e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6750 $Y=0.0970 $X2=0.6750 $Y2=0.1075
r60 26 47 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0970 $X2=0.6750 $Y2=0.0880
r61 44 45 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1205 $X2=0.6750 $Y2=0.1330
r62 43 44 0.867186 $w=1.3625e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.6750 $Y=0.1165 $X2=0.6750 $Y2=0.1205
r63 32 43 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1075 $X2=0.6750 $Y2=0.1165
r64 42 43 6.81353 $w=1.30847e-08 $l=3.89391e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7130 $Y=0.1080 $X2=0.6750 $Y2=0.1165
r65 41 42 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.7445
+ $Y=0.1080 $X2=0.7130 $Y2=0.1080
r66 40 41 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.1080 $X2=0.7445 $Y2=0.1080
r67 27 38 8.26388 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7965 $Y=0.1080 $X2=0.8370 $Y2=0.1080
r68 27 40 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.7965
+ $Y=0.1080 $X2=0.7560 $Y2=0.1080
r69 33 37 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1205 $X2=0.8370 $Y2=0.1330
r70 33 38 1.73456 $w=1.66e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8370 $Y=0.1205 $X2=0.8370 $Y2=0.1080
r71 15 3 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.8370
+ $Y=0.1350 $X2=0.8370 $Y2=0.1350
r72 3 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8370 $Y=0.1350
+ $X2=0.8370 $Y2=0.1330
.ends


*
.SUBCKT ICGx2_ASAP7_75t_R VSS VDD ENA SE CLK GCLK
*
* VSS VSS
* VDD VDD
* ENA ENA
* SE SE
* CLK CLK
* GCLK GCLK
*
*

MM19 N_MM19_d N_MM19_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM27 N_MM27_d N_MM18_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM10_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM6 N_MM6_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM20 N_MM20_d N_MM21_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM12 N_MM12_d N_MM0_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM13 N_MM13_d N_MM16_g N_MM13_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM14 N_MM14_d N_MM14_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24 N_MM24_d N_MM24_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@2 N_MM24@2_d N_MM24@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM26 N_MM26_d N_MM19_g N_MM26_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM18 N_MM18_d N_MM18_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM21 N_MM21_d N_MM21_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM16 N_MM16_d N_MM16_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM16@2 N_MM16@2_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM0@2 N_MM0@2_d N_MM14_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM25 N_MM25_d N_MM24_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@2 N_MM25@2_d N_MM24@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "ICGx2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "ICGx2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_ICGx2_ASAP7_75t_R%NOS1 VSS N_MM26_s N_MM18_d N_NOS1_1
+ PM_ICGx2_ASAP7_75t_R%NOS1
cc_1 N_NOS1_1 N_MM19_g 0.0125292f
cc_2 N_NOS1_1 N_MM18_g 0.0125758f
x_PM_ICGx2_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_ICGx2_ASAP7_75t_R%noxref_19
cc_3 N_noxref_19_1 N_MM19_g 0.00393361f
cc_4 N_noxref_19_1 N_NET0121_10 0.000401679f
x_PM_ICGx2_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_ICGx2_ASAP7_75t_R%noxref_20
cc_5 N_noxref_20_1 N_MM19_g 0.00393331f
cc_6 N_noxref_20_1 N_NET0121_11 0.0276625f
cc_7 N_noxref_20_1 N_noxref_19_1 0.00208735f
x_PM_ICGx2_ASAP7_75t_R%SE VSS SE N_MM18_g N_SE_1 N_SE_4 PM_ICGx2_ASAP7_75t_R%SE
cc_8 N_SE_1 N_ENA_1 0.00169567f
cc_9 N_SE_4 N_ENA_4 0.00520391f
cc_10 N_MM18_g N_MM19_g 0.00985307f
x_PM_ICGx2_ASAP7_75t_R%ENA VSS ENA N_MM19_g N_ENA_1 N_ENA_4
+ PM_ICGx2_ASAP7_75t_R%ENA
x_PM_ICGx2_ASAP7_75t_R%noxref_26 VSS N_noxref_26_1
+ PM_ICGx2_ASAP7_75t_R%noxref_26
cc_11 N_noxref_26_1 N_MM24@2_g 0.00146154f
cc_12 N_noxref_26_1 N_GCLK_8 0.000838657f
cc_13 N_noxref_26_1 N_noxref_25_1 0.00177248f
x_PM_ICGx2_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_ICGx2_ASAP7_75t_R%noxref_25
cc_14 N_noxref_25_1 N_MM24@2_g 0.00146165f
cc_15 N_noxref_25_1 N_GCLK_7 0.000841675f
x_PM_ICGx2_ASAP7_75t_R%GCLK VSS GCLK N_MM24_d N_MM24@2_d N_MM25_d N_MM25@2_d
+ N_GCLK_7 N_GCLK_8 N_GCLK_11 N_GCLK_1 N_GCLK_2 N_GCLK_10 N_GCLK_9
+ PM_ICGx2_ASAP7_75t_R%GCLK
cc_16 N_GCLK_7 N_GCLKN_18 0.000856101f
cc_17 N_GCLK_8 N_MM24@2_g 0.0309889f
cc_18 N_GCLK_11 N_GCLKN_1 0.00112187f
cc_19 N_GCLK_1 N_GCLKN_20 0.00179976f
cc_20 N_GCLK_1 N_MM24@2_g 0.00230692f
cc_21 N_GCLK_2 N_MM24@2_g 0.00237981f
cc_22 N_GCLK_10 N_GCLKN_23 0.00249155f
cc_23 N_GCLK_9 N_GCLKN_22 0.00305009f
cc_24 N_GCLK_8 N_GCLKN_1 0.00458536f
cc_25 N_GCLK_7 N_MM24_g 0.0372287f
cc_26 N_GCLK_7 N_MM24@2_g 0.0698178f
x_PM_ICGx2_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_ICGx2_ASAP7_75t_R%noxref_21
cc_27 N_noxref_21_1 N_CLKN_10 0.000837518f
cc_28 N_noxref_21_1 N_MS_3 0.00100914f
cc_29 N_noxref_21_1 N_MS_10 0.0169534f
cc_30 N_noxref_21_1 N_MM7_g 0.00534818f
x_PM_ICGx2_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_ICGx2_ASAP7_75t_R%noxref_22
cc_31 N_noxref_22_1 N_CLKN_11 0.000956656f
cc_32 N_noxref_22_1 N_MS_11 0.0170564f
cc_33 N_noxref_22_1 N_MM7_g 0.00577904f
cc_34 N_noxref_22_1 N_noxref_21_1 0.00153657f
x_PM_ICGx2_ASAP7_75t_R%NET0121 VSS N_MM3_g N_MM19_d N_MM27_d N_MM26_d
+ N_NET0121_11 N_NET0121_13 N_NET0121_4 N_NET0121_3 N_NET0121_12 N_NET0121_10
+ N_NET0121_1 N_NET0121_14 PM_ICGx2_ASAP7_75t_R%NET0121
cc_35 N_NET0121_11 N_ENA_1 0.000579346f
cc_36 N_NET0121_13 N_ENA_4 0.000668576f
cc_37 N_NET0121_4 N_MM19_g 0.000750777f
cc_38 N_NET0121_3 N_MM19_g 0.00108943f
cc_39 N_NET0121_12 N_ENA_4 0.0014352f
cc_40 N_NET0121_4 N_ENA_4 0.00303861f
cc_41 N_NET0121_11 N_MM19_g 0.0111053f
cc_42 N_NET0121_10 N_MM19_g 0.0403051f
cc_43 N_NET0121_1 N_MM18_g 0.00097167f
cc_44 N_NET0121_13 N_SE_4 0.00102799f
cc_45 N_NET0121_1 N_SE_1 0.00119135f
cc_46 N_NET0121_12 N_SE_4 0.0012138f
cc_47 N_NET0121_10 N_MM18_g 0.0109236f
cc_48 N_NET0121_14 N_SE_4 0.00753963f
cc_49 N_MM3_g N_MM18_g 0.0186749f
x_PM_ICGx2_ASAP7_75t_R%PU1 VSS N_MM3_d N_MM1_s N_PU1_3 N_PU1_1
+ PM_ICGx2_ASAP7_75t_R%PU1
cc_50 N_PU1_3 N_NET0121_1 0.000627824f
cc_51 N_PU1_3 N_MM3_g 0.0348994f
cc_52 N_PU1_3 N_CLK_15 0.000334704f
cc_53 N_PU1_3 N_CLK_1 0.000513634f
cc_54 N_PU1_3 N_MM1_g 0.0336043f
cc_55 N_PU1_1 N_MH_18 0.00109775f
cc_56 N_PU1_1 N_MH_7 0.00288966f
x_PM_ICGx2_ASAP7_75t_R%PD3 VSS N_MM9_s N_MM8_d N_PD3_3 N_PD3_1
+ PM_ICGx2_ASAP7_75t_R%PD3
cc_57 N_PD3_3 N_MM9_g 0.0146719f
cc_58 N_PD3_3 N_MM11_g 0.0162355f
cc_59 N_PD3_1 N_MH_22 0.000207234f
cc_60 N_PD3_1 N_MH_16 0.00061144f
cc_61 N_PD3_1 N_MH_24 0.000307959f
cc_62 N_PD3_1 N_MH_8 0.00212167f
x_PM_ICGx2_ASAP7_75t_R%NET0140 VSS N_MM2_s N_MM14_d N_NET0140_1
+ PM_ICGx2_ASAP7_75t_R%NET0140
cc_63 N_NET0140_1 N_MM2_g 0.0173194f
cc_64 N_NET0140_1 N_MM14_g 0.0173193f
x_PM_ICGx2_ASAP7_75t_R%PD1 VSS N_MM5_d N_MM4_s N_PD1_4 N_PD1_5 N_PD1_1
+ PM_ICGx2_ASAP7_75t_R%PD1
cc_65 N_PD1_4 N_NET0121_1 0.000768702f
cc_66 N_PD1_4 N_MM3_g 0.0359384f
cc_67 N_PD1_5 N_CLK_1 0.00231372f
cc_68 N_PD1_5 N_MM1_g 0.0732003f
cc_69 N_PD1_5 N_CLKN_1 0.000683195f
cc_70 N_PD1_5 N_CLKN_14 0.00272143f
cc_71 N_PD1_5 N_MM10_g 0.0334571f
cc_72 N_PD1_1 N_MH_8 0.00133112f
cc_73 N_PD1_1 N_MH_16 0.0029334f
x_PM_ICGx2_ASAP7_75t_R%NET0141 VSS N_MM12_d N_MM13_s N_NET0141_1
+ PM_ICGx2_ASAP7_75t_R%NET0141
cc_74 N_NET0141_1 N_MM16_g 0.0174349f
cc_75 N_NET0141_1 N_MM0_g 0.0172741f
x_PM_ICGx2_ASAP7_75t_R%PD2 VSS N_MM10_s N_MM11_d N_PD2_5 N_PD2_4 N_PD2_1
+ PM_ICGx2_ASAP7_75t_R%PD2
cc_76 N_PD2_5 N_CLK_8 0.000220944f
cc_77 N_PD2_4 N_MM9_g 0.00732298f
cc_78 N_PD2_1 N_MM9_g 0.000993903f
cc_79 N_PD2_5 N_MM9_g 0.0237224f
cc_80 N_PD2_1 N_MM10_g 0.000492672f
cc_81 N_PD2_4 N_MM10_g 0.0149721f
cc_82 N_PD2_5 N_MM11_g 0.0149322f
cc_83 N_PD2_1 N_MH_22 9.5354e-20
cc_84 N_PD2_1 N_MH_7 0.000117211f
cc_85 N_PD2_1 N_MH_23 0.000256153f
cc_86 N_PD2_1 N_MH_25 0.000296432f
cc_87 N_PD2_4 N_MH_18 0.000643007f
cc_88 N_PD2_1 N_MH_20 0.000491752f
cc_89 N_PD2_4 N_MH_7 0.000618538f
cc_90 N_PD2_1 N_MH_30 0.002704f
x_PM_ICGx2_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_ICGx2_ASAP7_75t_R%noxref_23
cc_91 N_noxref_23_1 N_MM21_g 0.00136326f
cc_92 N_noxref_23_1 N_CLKN_10 0.0376459f
cc_93 N_noxref_23_1 N_MS_10 0.000573045f
cc_94 N_noxref_23_1 N_noxref_21_1 0.00773065f
cc_95 N_noxref_23_1 N_noxref_22_1 0.000477264f
x_PM_ICGx2_ASAP7_75t_R%GCLKN VSS N_MM24_g N_MM24@2_g N_MM2_d N_MM13_d
+ N_MM16@2_d N_MM0@2_d N_MM0_d N_MM16_d N_GCLKN_14 N_GCLKN_5 N_GCLKN_15
+ N_GCLKN_3 N_GCLKN_17 N_GCLKN_4 N_GCLKN_16 N_GCLKN_18 N_GCLKN_21 N_GCLKN_1
+ N_GCLKN_20 N_GCLKN_23 N_GCLKN_22 PM_ICGx2_ASAP7_75t_R%GCLKN
cc_96 N_GCLKN_14 N_CLK_22 0.000418721f
cc_97 N_GCLKN_14 N_CLK_23 0.000181372f
cc_98 N_GCLKN_14 N_CLK_18 0.000292382f
cc_99 N_GCLKN_5 N_CLK_4 0.000341215f
cc_100 N_GCLKN_15 N_MM16_g 0.011547f
cc_101 N_GCLKN_3 N_CLK_17 0.000420541f
cc_102 N_GCLKN_17 N_CLK_18 0.000484965f
cc_103 N_GCLKN_5 N_MM2_g 0.00088628f
cc_104 N_GCLKN_3 N_MM16_g 0.00126558f
cc_105 N_GCLKN_4 N_MM2_g 0.00150636f
cc_106 N_GCLKN_16 N_CLK_4 0.00246685f
cc_107 N_GCLKN_17 N_CLK_17 0.00259149f
cc_108 N_GCLKN_17 N_CLK_22 0.00384972f
cc_109 N_GCLKN_16 N_MM2_g 0.0109938f
cc_110 N_GCLKN_14 N_MM16_g 0.0332745f
cc_111 N_GCLKN_14 N_MM2_g 0.0657895f
cc_112 N_GCLKN_15 N_MH_32 0.00011382f
cc_113 N_GCLKN_15 N_MH_2 0.000447009f
cc_114 N_GCLKN_15 N_MH_31 0.000154528f
cc_115 N_GCLKN_15 N_MH_33 0.000496051f
cc_116 N_GCLKN_14 N_MM14_g 0.00030072f
cc_117 N_GCLKN_16 N_MM14_g 0.0112374f
cc_118 N_GCLKN_18 N_MH_26 0.00037162f
cc_119 N_GCLKN_5 N_MM14_g 0.000402063f
cc_120 N_GCLKN_3 N_MM0_g 0.000411282f
cc_121 N_GCLKN_21 N_MH_33 0.000496759f
cc_122 N_GCLKN_4 N_MH_27 0.00182649f
cc_123 N_GCLKN_1 N_MH_3 0.00250238f
cc_124 N_GCLKN_18 N_MH_33 0.00135518f
cc_125 N_GCLKN_20 N_MH_33 0.00270788f
cc_126 N_GCLKN_18 N_MH_27 0.00990882f
cc_127 N_MM24_g N_MM14_g 0.0172029f
cc_128 N_GCLKN_15 N_MM0_g 0.0253868f
x_PM_ICGx2_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_ICGx2_ASAP7_75t_R%noxref_24
cc_129 N_noxref_24_1 N_MM21_g 0.00136824f
cc_130 N_noxref_24_1 N_CLKN_4 0.00041051f
cc_131 N_noxref_24_1 N_CLKN_11 0.0373735f
cc_132 N_noxref_24_1 N_MS_11 0.000538368f
cc_133 N_noxref_24_1 N_noxref_21_1 0.000473227f
cc_134 N_noxref_24_1 N_noxref_22_1 0.00777077f
cc_135 N_noxref_24_1 N_noxref_23_1 0.00123136f
x_PM_ICGx2_ASAP7_75t_R%CLK VSS CLK N_MM1_g N_MM9_g N_MM21_g N_MM16_g N_MM2_g
+ N_CLK_23 N_CLK_1 N_CLK_15 N_CLK_21 N_CLK_20 N_CLK_16 N_CLK_8 N_CLK_17 N_CLK_3
+ N_CLK_2 N_CLK_19 N_CLK_22 N_CLK_4 N_CLK_18 PM_ICGx2_ASAP7_75t_R%CLK
cc_136 N_CLK_23 N_NET0121_14 0.000640938f
cc_137 N_CLK_1 N_NET0121_1 0.00159338f
cc_138 N_MM1_g N_MM3_g 0.00327231f
cc_139 N_CLK_15 N_NET0121_14 0.00460273f
x_PM_ICGx2_ASAP7_75t_R%MS VSS N_MM11_g N_MM6_d N_MM7_d N_MS_1 N_MS_12 N_MS_13
+ N_MS_15 N_MS_3 N_MS_14 N_MS_4 N_MS_11 N_MS_10 PM_ICGx2_ASAP7_75t_R%MS
cc_140 N_MM11_g N_CLK_20 0.000217535f
cc_141 N_MM11_g N_CLK_23 0.000125382f
cc_142 N_MM11_g N_CLK_8 0.00294032f
cc_143 N_MS_1 N_CLK_19 0.000552116f
cc_144 N_MS_1 N_CLK_8 0.00153715f
cc_145 N_MS_12 N_CLK_20 0.000626225f
cc_146 N_MS_13 N_CLK_23 0.00150955f
cc_147 N_MS_12 N_CLK_23 0.00158104f
cc_148 N_MS_12 N_CLK_19 0.00255784f
cc_149 N_MM11_g N_MM9_g 0.0131881f
cc_150 N_MS_13 N_CLKN_11 0.000122571f
cc_151 N_MS_13 N_CLKN_16 0.000223071f
cc_152 N_MS_15 N_CLKN_3 0.00024744f
cc_153 N_MS_3 N_CLKN_16 0.000253119f
cc_154 N_MS_13 N_CLKN_4 0.000275436f
cc_155 N_MS_14 N_CLKN_17 0.000855618f
cc_156 N_MS_15 N_CLKN_16 0.000951897f
cc_157 N_MS_14 N_CLKN_18 0.00147397f
cc_158 N_MS_13 N_CLKN_13 0.00669086f
x_PM_ICGx2_ASAP7_75t_R%CLKN VSS N_MM10_g N_MM20_d N_MM21_d N_CLKN_10 N_CLKN_13
+ N_CLKN_18 N_CLKN_3 N_CLKN_15 N_CLKN_12 N_CLKN_1 N_CLKN_17 N_CLKN_11 N_CLKN_14
+ N_CLKN_16 N_CLKN_4 PM_ICGx2_ASAP7_75t_R%CLKN
cc_159 N_CLKN_10 N_CLK_21 0.000185119f
cc_160 N_CLKN_13 N_CLK_21 0.000185189f
cc_161 N_CLKN_18 N_CLK_20 0.000263922f
cc_162 N_CLKN_3 N_CLK_16 0.000285932f
cc_163 N_CLKN_15 N_CLK_15 0.000293691f
cc_164 N_CLKN_12 N_CLK_15 0.00409448f
cc_165 N_CLKN_1 N_CLK_8 0.000315533f
cc_166 N_CLKN_13 N_CLK_16 0.00501322f
cc_167 N_CLKN_1 N_CLK_1 0.0015249f
cc_168 N_CLKN_17 N_CLK_17 0.000464453f
cc_169 N_CLKN_11 N_MM21_g 0.0157643f
cc_170 N_CLKN_15 N_CLK_23 0.000516958f
cc_171 N_CLKN_13 N_CLK_23 0.000698225f
cc_172 N_CLKN_14 N_CLK_15 0.000812026f
cc_173 N_CLKN_16 N_CLK_16 0.00093557f
cc_174 N_CLKN_3 N_MM21_g 0.00094502f
cc_175 N_CLKN_3 N_CLK_3 0.000965282f
cc_176 N_CLKN_4 N_MM21_g 0.00135352f
cc_177 N_CLKN_1 N_CLK_2 0.00147977f
cc_178 N_MM10_g N_MM1_g 0.00161597f
cc_179 N_CLKN_11 N_CLK_3 0.0016435f
cc_180 N_CLKN_17 N_CLK_21 0.00174329f
cc_181 N_MM10_g N_MM9_g 0.00910327f
cc_182 N_CLKN_18 N_CLK_23 0.0259678f
cc_183 N_CLKN_10 N_MM21_g 0.0541723f
x_PM_ICGx2_ASAP7_75t_R%MH VSS N_MM7_g N_MM0_g N_MM14_g N_MM4_d N_MM9_d N_MM1_d
+ N_MM10_d N_MH_23 N_MH_7 N_MH_21 N_MH_29 N_MH_19 N_MH_17 N_MH_27 N_MH_32
+ N_MH_33 N_MH_18 N_MH_3 N_MH_1 N_MH_25 N_MH_26 N_MH_20 N_MH_22 N_MH_24 N_MH_16
+ N_MH_8 N_MH_2 N_MH_30 N_MH_31 PM_ICGx2_ASAP7_75t_R%MH
cc_184 N_MH_23 N_CLK_19 7.89505e-20
cc_185 N_MH_7 N_CLK_15 0.00084019f
cc_186 N_MH_21 N_MM9_g 0.000133524f
cc_187 N_MH_29 N_CLK_19 0.000143071f
cc_188 N_MH_19 N_MM1_g 0.00014953f
cc_189 N_MH_17 N_MM9_g 0.000175721f
cc_190 N_MH_27 N_CLK_22 0.000201848f
cc_191 N_MH_7 N_CLK_1 0.000204324f
cc_192 N_MH_32 N_CLK_16 0.00305637f
cc_193 N_MH_33 N_CLK_4 0.00024448f
cc_194 N_MH_18 N_MM1_g 0.0338856f
cc_195 N_MH_3 N_CLK_4 0.000264041f
cc_196 N_MH_1 N_CLK_8 0.000271258f
cc_197 N_MH_1 N_CLK_20 0.000305803f
cc_198 N_MH_25 N_CLK_20 0.00476149f
cc_199 N_MH_26 N_CLK_16 0.000362305f
cc_200 N_MH_27 N_CLK_4 0.000401496f
cc_201 N_MH_20 N_CLK_15 0.000487324f
cc_202 N_MH_22 N_CLK_8 0.00250082f
cc_203 N_MM7_g N_CLK_8 0.00054433f
cc_204 N_MH_3 N_MM2_g 0.000562701f
cc_205 N_MH_18 N_CLK_1 0.000569951f
cc_206 N_MH_24 N_CLK_23 0.000708792f
cc_207 N_MH_16 N_CLK_2 0.000886988f
cc_208 N_MH_8 N_MM9_g 0.00101642f
cc_209 N_MH_7 N_MM1_g 0.0011796f
cc_210 N_MH_2 N_CLK_3 0.00305765f
cc_211 N_MH_25 N_CLK_19 0.00140162f
cc_212 N_MH_32 N_CLK_17 0.00148925f
cc_213 N_MM14_g N_CLK_4 0.00166613f
cc_214 N_MM0_g N_MM21_g 0.00166641f
cc_215 N_MH_25 N_CLK_23 0.00236986f
cc_216 N_MH_22 N_CLK_19 0.00383142f
cc_217 N_MH_27 N_CLK_18 0.00388213f
cc_218 N_MM14_g N_MM2_g 0.0071603f
cc_219 N_MM0_g N_MM16_g 0.00886723f
cc_220 N_MH_16 N_MM9_g 0.0366414f
cc_221 N_MM0_g N_MM10_g 0.000126632f
cc_222 N_MH_27 N_MM10_g 8.92997e-20
cc_223 N_MM7_g N_MM10_g 9.38751e-20
cc_224 N_MH_17 N_MM10_g 0.000144983f
cc_225 N_MH_32 N_CLKN_16 0.000149975f
cc_226 N_MH_19 N_MM10_g 0.000166264f
cc_227 N_MH_8 N_CLKN_14 0.000186868f
cc_228 N_MH_7 N_CLKN_15 0.000193659f
cc_229 N_MH_30 N_CLKN_15 0.000197599f
cc_230 N_MH_26 N_CLKN_16 0.000214968f
cc_231 N_MH_25 N_CLKN_13 0.000249005f
cc_232 N_MH_24 N_CLKN_3 0.00111962f
cc_233 N_MH_18 N_MM10_g 0.0166804f
cc_234 N_MH_20 N_CLKN_15 0.00477988f
cc_235 N_MH_23 N_CLKN_15 0.000541385f
cc_236 N_MH_29 N_CLKN_15 0.000688789f
cc_237 N_MH_8 N_CLKN_1 0.000701545f
cc_238 N_MH_8 N_MM10_g 0.00133706f
cc_239 N_MH_7 N_MM10_g 0.00142321f
cc_240 N_MH_16 N_CLKN_1 0.00148257f
cc_241 N_MH_21 N_CLKN_14 0.00191012f
cc_242 N_MH_25 N_CLKN_18 0.00329975f
cc_243 N_MH_22 N_CLKN_12 0.00379313f
cc_244 N_MH_24 N_CLKN_16 0.00436117f
cc_245 N_MH_16 N_MM10_g 0.0536179f
cc_246 N_MH_8 N_MM11_g 0.000202446f
cc_247 N_MH_24 N_MM11_g 0.000315363f
cc_248 N_MH_1 N_MS_4 0.00197807f
cc_249 N_MM7_g N_MS_1 0.000552093f
cc_250 N_MH_24 N_MS_1 0.000727436f
cc_251 N_MH_1 N_MS_11 0.0012631f
cc_252 N_MH_22 N_MS_12 0.00130815f
cc_253 N_MH_25 N_MS_13 0.0013873f
cc_254 N_MM7_g N_MS_3 0.00170061f
cc_255 N_MH_25 N_MS_14 0.00239907f
cc_256 N_MM7_g N_MS_10 0.00643105f
cc_257 N_MM7_g N_MS_11 0.00675895f
cc_258 N_MH_24 N_MS_12 0.0036925f
cc_259 N_MH_24 N_MS_15 0.00539924f
cc_260 N_MM7_g N_MM11_g 0.0297137f
*END of ICGx2_ASAP7_75t_R.pxi
.ENDS
** Design:	ICGx3_ASAP7_75t_R
* Created:	"Fri Aug 17 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "ICGx3_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "ICGx3_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_ICGx3_ASAP7_75t_R%NOS1 VSS 2 3 1
c1 1 VSS 0.00087961f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2160 $X2=0.1080 $Y2=0.2160
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2160 $X2=0.1080 $Y2=0.2160
.ends

.subckt PM_ICGx3_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.0320326f
.ends

.subckt PM_ICGx3_ASAP7_75t_R%ENA VSS 8 3 1 4
c1 1 VSS 0.00207589f
c2 3 VSS 0.0329499f
c3 4 VSS 0.00973895f
r1 9 10 2.3902 $w=1.3e-08 $l=1.03e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1267 $X2=0.0810 $Y2=0.1370
r2 8 9 0.408082 $w=1.3e-08 $l=1.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1250 $X2=0.0810 $Y2=0.1267
r3 8 4 6.47102 $w=1.3e-08 $l=2.78e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1250 $X2=0.0810 $Y2=0.0972
r4 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r5 1 10 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1370
.ends

.subckt PM_ICGx3_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.00478249f
.ends

.subckt PM_ICGx3_ASAP7_75t_R%SE VSS 8 3 1 4
c1 1 VSS 0.00634763f
c2 3 VSS 0.0830419f
c3 4 VSS 0.00452691f
r1 9 10 2.3902 $w=1.3e-08 $l=1.03e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1267 $X2=0.1350 $Y2=0.1370
r2 8 9 0.408082 $w=1.3e-08 $l=1.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1250 $X2=0.1350 $Y2=0.1267
r3 8 4 6.47102 $w=1.3e-08 $l=2.78e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1250 $X2=0.1350 $Y2=0.0972
r4 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r5 1 10 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1370
.ends

.subckt PM_ICGx3_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.00532282f
.ends

.subckt PM_ICGx3_ASAP7_75t_R%noxref_26 VSS 1
c1 1 VSS 0.0056434f
.ends

.subckt PM_ICGx3_ASAP7_75t_R%GCLK VSS 32 24 25 36 44 45 47 13 17 3 15 4 1 2 18
+ 16 14
c1 1 VSS 0.00990947f
c2 2 VSS 0.00992067f
c3 3 VSS 0.00798639f
c4 4 VSS 0.00797052f
c5 13 VSS 0.00459114f
c6 14 VSS 0.00348501f
c7 15 VSS 0.0045078f
c8 16 VSS 0.00343086f
c9 17 VSS 0.0166448f
c10 18 VSS 0.0140382f
c11 19 VSS 0.00359745f
c12 20 VSS 0.00281678f
c13 21 VSS 0.00286572f
r1 16 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0115 $Y=0.2025 $X2=1.0240 $Y2=0.2025
r2 47 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0090 $Y=0.2025 $X2=1.0115 $Y2=0.2025
r3 45 43 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9350 $Y=0.2025 $X2=0.9325 $Y2=0.2025
r4 2 43 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9180 $Y=0.2025 $X2=0.9325 $Y2=0.2025
r5 15 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9035 $Y=0.2025 $X2=0.9180 $Y2=0.2025
r6 44 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9010 $Y=0.2025 $X2=0.9035 $Y2=0.2025
r7 4 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0260 $Y=0.2025
+ $X2=1.0260 $Y2=0.2340
r8 2 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.9180 $Y=0.2025
+ $X2=0.9180 $Y2=0.2340
r9 39 40 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.2340 $X2=1.0395 $Y2=0.2340
r10 38 39 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.9720
+ $Y=0.2340 $X2=1.0260 $Y2=0.2340
r11 37 38 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.2340 $X2=0.9720 $Y2=0.2340
r12 18 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.9045
+ $Y=0.2340 $X2=0.9180 $Y2=0.2340
r13 21 34 2.6649 $w=1.77676e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0530 $Y=0.2340 $X2=1.0530 $Y2=0.2155
r14 21 40 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0530 $Y=0.2340 $X2=1.0395 $Y2=0.2340
r15 14 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.0115 $Y=0.0675 $X2=1.0240 $Y2=0.0675
r16 36 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.0090 $Y=0.0675 $X2=1.0115 $Y2=0.0675
r17 33 34 6.8208 $w=1.3e-08 $l=2.93e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1862 $X2=1.0530 $Y2=0.2155
r18 32 33 4.72209 $w=1.3e-08 $l=2.02e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1660 $X2=1.0530 $Y2=0.1862
r19 32 31 12.0676 $w=1.3e-08 $l=5.18e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1660 $X2=1.0530 $Y2=0.1142
r20 19 20 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.0540 $X2=1.0530 $Y2=0.0360
r21 19 31 14.0497 $w=1.3e-08 $l=6.02e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.0540 $X2=1.0530 $Y2=0.1142
r22 3 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0260 $Y=0.0675
+ $X2=1.0260 $Y2=0.0360
r23 20 30 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0530 $Y=0.0360 $X2=1.0395 $Y2=0.0360
r24 29 30 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.0360 $X2=1.0395 $Y2=0.0360
r25 28 29 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.9720
+ $Y=0.0360 $X2=1.0260 $Y2=0.0360
r26 27 28 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.0360 $X2=0.9720 $Y2=0.0360
r27 26 27 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.9045
+ $Y=0.0360 $X2=0.9180 $Y2=0.0360
r28 17 26 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.8895
+ $Y=0.0360 $X2=0.9045 $Y2=0.0360
r29 1 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.9180 $Y=0.0675
+ $X2=0.9180 $Y2=0.0360
r30 25 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9350 $Y=0.0675 $X2=0.9325 $Y2=0.0675
r31 1 23 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9180 $Y=0.0675 $X2=0.9325 $Y2=0.0675
r32 13 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9035 $Y=0.0675 $X2=0.9180 $Y2=0.0675
r33 24 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9010 $Y=0.0675 $X2=0.9035 $Y2=0.0675
.ends

.subckt PM_ICGx3_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.00364721f
.ends

.subckt PM_ICGx3_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.00366229f
.ends

.subckt PM_ICGx3_ASAP7_75t_R%NET056 VSS 2 3 1
c1 1 VSS 0.000863663f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.0675 $X2=0.7020 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.0675 $X2=0.7020 $Y2=0.0675
.ends

.subckt PM_ICGx3_ASAP7_75t_R%PD3 VSS 5 8 3 1
c1 1 VSS 0.00335282f
c2 3 VSS 0.00246954f
r1 8 7 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0405 $X2=0.3925 $Y2=0.0405
r2 1 7 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3800 $Y=0.0405 $X2=0.3925 $Y2=0.0405
r3 4 1 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3680 $Y=0.0405 $X2=0.3800 $Y2=0.0405
r4 3 4 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.0405 $X2=0.3680 $Y2=0.0405
r5 5 3 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0405 $X2=0.3635 $Y2=0.0405
.ends

.subckt PM_ICGx3_ASAP7_75t_R%PU1 VSS 5 8 3 1
c1 1 VSS 0.00536713f
c2 3 VSS 0.00340052f
r1 8 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r2 6 7 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2260 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r3 1 6 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2140 $Y=0.2025 $X2=0.2260 $Y2=0.2025
r4 3 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2140 $Y2=0.2025
r5 5 3 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
.ends

.subckt PM_ICGx3_ASAP7_75t_R%MS VSS 9 40 46 1 12 13 15 3 14 4 11 10
c1 1 VSS 0.00206478f
c2 3 VSS 0.00502444f
c3 4 VSS 0.0060284f
c4 9 VSS 0.0369145f
c5 10 VSS 0.00304752f
c6 11 VSS 0.00308632f
c7 12 VSS 0.00122221f
c8 13 VSS 0.00123971f
c9 14 VSS 0.00665295f
c10 15 VSS 0.000343258f
r1 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2295 $X2=0.4840 $Y2=0.2295
r2 46 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2295 $X2=0.4715 $Y2=0.2295
r3 4 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2295
+ $X2=0.4860 $Y2=0.2330
r4 42 43 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.2330 $X2=0.4990 $Y2=0.2330
r5 14 38 1.06916 $w=1.78e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.2330 $X2=0.5125 $Y2=0.2235
r6 14 43 1.90218 $w=1.65185e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5125 $Y=0.2330 $X2=0.4990 $Y2=0.2330
r7 10 31 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0405 $X2=0.4840 $Y2=0.0405
r8 40 10 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0405 $X2=0.4715 $Y2=0.0405
r9 37 38 2.49333 $w=1.4e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.2110 $X2=0.5125 $Y2=0.2235
r10 36 37 4.1888 $w=1.4e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.1900 $X2=0.5125 $Y2=0.2110
r11 35 36 3.69013 $w=1.4e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.1715 $X2=0.5125 $Y2=0.1900
r12 34 35 3.69013 $w=1.4e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.1530 $X2=0.5125 $Y2=0.1715
r13 33 34 4.1888 $w=1.4e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.1320 $X2=0.5125 $Y2=0.1530
r14 32 33 4.88693 $w=1.4e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.1075 $X2=0.5125 $Y2=0.1320
r15 13 15 0.843012 $w=1.80909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5125 $Y=0.0930 $X2=0.5125 $Y2=0.0820
r16 13 32 2.89227 $w=1.4e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.0930 $X2=0.5125 $Y2=0.1075
r17 3 29 10.904 $w=2.02e-08 $l=1.85e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4860 $Y=0.0635 $X2=0.4860 $Y2=0.0820
r18 3 31 13.5563 $w=2.02e-08 $l=2.3e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4860 $Y=0.0635 $X2=0.4860 $Y2=0.0405
r19 15 28 1.37684 $w=2.03185e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5125 $Y=0.0820 $X2=0.4990 $Y2=0.0820
r20 27 28 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.0820 $X2=0.4990 $Y2=0.0820
r21 27 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0820
+ $X2=0.4860 $Y2=0.0820
r22 26 27 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4750
+ $Y=0.0820 $X2=0.4860 $Y2=0.0820
r23 25 26 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4600
+ $Y=0.0820 $X2=0.4750 $Y2=0.0820
r24 24 25 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4310
+ $Y=0.0820 $X2=0.4600 $Y2=0.0820
r25 23 24 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.4145
+ $Y=0.0820 $X2=0.4310 $Y2=0.0820
r26 21 23 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4055
+ $Y=0.0820 $X2=0.4145 $Y2=0.0820
r27 12 21 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3965
+ $Y=0.0820 $X2=0.4055 $Y2=0.0820
r28 18 20 2.94116 $w=2.133e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.4060
+ $Y=0.0820 $X2=0.4160 $Y2=0.0820
r29 18 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4060 $Y=0.0820
+ $X2=0.4055 $Y2=0.0820
r30 1 18 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.3960
+ $Y=0.0820 $X2=0.4060 $Y2=0.0820
r31 1 19 0.851883 $w=1.865e-08 $l=2e-09 $layer=LIG $thickness=4.8e-08 $X=0.3960
+ $Y=0.0820 $X2=0.3940 $Y2=0.0820
r32 17 18 2.35044 $w=2.2e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.4050
+ $Y=0.0820 $X2=0.4060 $Y2=0.0820
r33 17 19 0.590723 $w=1.53e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4050 $Y=0.0820 $X2=0.3940 $Y2=0.0820
r34 17 20 0.590723 $w=1.53e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4050 $Y=0.0820 $X2=0.4160 $Y2=0.0820
r35 9 17 0.314665 $w=2.27e-07 $l=5.3e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4050 $Y2=0.0820
.ends

.subckt PM_ICGx3_ASAP7_75t_R%PD1 VSS 7 10 4 5 1
c1 1 VSS 0.00979402f
c2 4 VSS 0.00323881f
c3 5 VSS 0.00185978f
r1 10 9 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r2 8 9 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2800 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r3 5 8 0.123457 $w=8.1e-08 $l=1e-08 $layer=N_src_drn $thickness=1e-09 $X=0.2700
+ $Y=0.0675 $X2=0.2800 $Y2=0.0675
r4 4 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0675 $X2=0.2140 $Y2=0.0675
r5 7 4 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2015 $Y2=0.0675
r6 1 5 1e-05
.ends

.subckt PM_ICGx3_ASAP7_75t_R%NET059 VSS 2 3 1
c1 1 VSS 0.000931854f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.0675 $X2=0.8100 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8270 $Y=0.0675 $X2=0.8100 $Y2=0.0675
.ends

.subckt PM_ICGx3_ASAP7_75t_R%PD2 VSS 7 13 5 4 1
c1 1 VSS 0.0072931f
c2 4 VSS 0.00188002f
c3 5 VSS 0.00238549f
r1 13 12 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r2 5 12 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3800 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r3 10 5 9.87715 $w=2.32e-08 $l=2.1e-08 $layer=LISD $thickness=2.7e-08 $X=0.3570
+ $Y=0.2295 $X2=0.3780 $Y2=0.2295
r4 9 10 6.11443 $w=2.32e-08 $l=1.3e-08 $layer=LISD $thickness=2.7e-08 $X=0.3440
+ $Y=0.2295 $X2=0.3570 $Y2=0.2295
r5 8 9 2.82204 $w=2.32e-08 $l=6e-09 $layer=LISD $thickness=2.7e-08 $X=0.3380
+ $Y=0.2295 $X2=0.3440 $Y2=0.2295
r6 1 8 6.58477 $w=2.32e-08 $l=1.4e-08 $layer=LISD $thickness=2.7e-08 $X=0.3240
+ $Y=0.2295 $X2=0.3380 $Y2=0.2295
r7 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2295 $X2=0.3220 $Y2=0.2295
r8 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2295 $X2=0.3095 $Y2=0.2295
.ends

.subckt PM_ICGx3_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.0042336f
.ends

.subckt PM_ICGx3_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.00441228f
.ends

.subckt PM_ICGx3_ASAP7_75t_R%MH VSS 13 14 15 77 81 100 104 23 7 21 29 19 17 27
+ 32 33 18 3 1 25 26 20 22 24 16 8 2 30 31
c1 1 VSS 0.0023512f
c2 2 VSS 0.0046007f
c3 3 VSS 0.00385685f
c4 7 VSS 0.00516563f
c5 8 VSS 0.00493236f
c6 13 VSS 0.036861f
c7 14 VSS 0.0818833f
c8 15 VSS 0.0817601f
c9 16 VSS 0.00317832f
c10 17 VSS 0.000556973f
c11 18 VSS 0.00315327f
c12 19 VSS 0.000592325f
c13 20 VSS 0.00828662f
c14 21 VSS 0.00485963f
c15 22 VSS 0.000832664f
c16 23 VSS 0.000426805f
c17 24 VSS 0.0293022f
c18 25 VSS 0.00200931f
c19 26 VSS 0.00222487f
c20 27 VSS 0.00201643f
c21 28 VSS 0.00226764f
c22 29 VSS 7.47383e-20
c23 30 VSS 0.00263428f
c24 31 VSS 0.00334412f
c25 32 VSS 0.000686684f
c26 33 VSS 0.00130036f
r1 104 103 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2295 $X2=0.2845 $Y2=0.2295
r2 102 103 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2800 $Y=0.2295 $X2=0.2845 $Y2=0.2295
r3 18 102 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2680 $Y=0.2295 $X2=0.2800 $Y2=0.2295
r4 19 18 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2295 $X2=0.2680 $Y2=0.2295
r5 98 99 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.1890 $X2=0.2600 $Y2=0.1890
r6 100 98 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.1890 $X2=0.2555 $Y2=0.1890
r7 18 99 0.185185 $w=5.4e-08 $l=1e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.1890 $X2=0.2600 $Y2=0.1890
r8 7 94 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2295
+ $X2=0.2700 $Y2=0.2320
r9 7 18 23.8708 $w=2.02e-08 $l=4.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.2700 $Y=0.2295 $X2=0.2700 $Y2=0.1890
r10 94 95 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2320 $X2=0.2835 $Y2=0.2320
r11 92 95 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3060
+ $Y=0.2320 $X2=0.2835 $Y2=0.2320
r12 20 30 2.96589 $w=1.31923e-08 $l=2.31193e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3365 $Y=0.2320 $X2=0.3580 $Y2=0.2235
r13 20 92 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.3365
+ $Y=0.2320 $X2=0.3060 $Y2=0.2320
r14 1 86 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1900
+ $X2=0.4590 $Y2=0.1900
r15 13 1 3.49039 $w=1.235e-07 $l=5.5e-08 $layer=LIG $thickness=5.2e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4590 $Y2=0.1900
r16 23 75 2.8493 $w=1.32e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.2110 $X2=0.3580 $Y2=0.1985
r17 23 30 2.8493 $w=1.32e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.2110 $X2=0.3580 $Y2=0.2235
r18 85 86 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4485
+ $Y=0.1900 $X2=0.4590 $Y2=0.1900
r19 84 85 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4305
+ $Y=0.1900 $X2=0.4485 $Y2=0.1900
r20 83 84 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1900 $X2=0.4305 $Y2=0.1900
r21 82 83 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3940
+ $Y=0.1900 $X2=0.4050 $Y2=0.1900
r22 25 29 3.78225 $w=1.50238e-08 $l=2.15058e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3795 $Y=0.1900 $X2=0.3580 $Y2=0.1895
r23 25 82 3.38125 $w=1.3e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3795
+ $Y=0.1900 $X2=0.3940 $Y2=0.1900
r24 81 80 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0405 $X2=0.3385 $Y2=0.0405
r25 79 80 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3340 $Y=0.0405 $X2=0.3385 $Y2=0.0405
r26 8 79 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3220 $Y=0.0405 $X2=0.3340 $Y2=0.0405
r27 17 8 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0405 $X2=0.3220 $Y2=0.0405
r28 16 8 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0810 $X2=0.3220 $Y2=0.0810
r29 77 16 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0810 $X2=0.3095 $Y2=0.0810
r30 29 70 0.983973 $w=1.77222e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.3580 $Y=0.1895 $X2=0.3580 $Y2=0.1805
r31 29 75 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.1895 $X2=0.3580 $Y2=0.1985
r32 8 63 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0405
+ $X2=0.3195 $Y2=0.0360
r33 69 70 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.1710 $X2=0.3580 $Y2=0.1805
r34 68 69 6.99569 $w=1.3e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.1410 $X2=0.3580 $Y2=0.1710
r35 67 68 8.27824 $w=1.3e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.1055 $X2=0.3580 $Y2=0.1410
r36 66 67 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.0905 $X2=0.3580 $Y2=0.1055
r37 65 66 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.0815 $X2=0.3580 $Y2=0.0905
r38 64 65 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.0725 $X2=0.3580 $Y2=0.0815
r39 22 28 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.0585 $X2=0.3580 $Y2=0.0360
r40 22 64 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.0585 $X2=0.3580 $Y2=0.0725
r41 21 61 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3285
+ $Y=0.0360 $X2=0.3410 $Y2=0.0360
r42 21 63 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3285
+ $Y=0.0360 $X2=0.3195 $Y2=0.0360
r43 28 60 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3580 $Y=0.0360 $X2=0.3795 $Y2=0.0360
r44 28 61 2.78392 $w=1.56471e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3580 $Y=0.0360 $X2=0.3410 $Y2=0.0360
r45 59 60 18.0722 $w=1.3e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.4570
+ $Y=0.0360 $X2=0.3795 $Y2=0.0360
r46 58 59 19.4713 $w=1.3e-08 $l=8.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5405
+ $Y=0.0360 $X2=0.4570 $Y2=0.0360
r47 57 58 10.1438 $w=1.3e-08 $l=4.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5840
+ $Y=0.0360 $X2=0.5405 $Y2=0.0360
r48 56 57 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.6105
+ $Y=0.0360 $X2=0.5840 $Y2=0.0360
r49 55 56 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0360 $X2=0.6105 $Y2=0.0360
r50 24 31 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6480 $Y=0.0360 $X2=0.6750 $Y2=0.0360
r51 24 55 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.6480
+ $Y=0.0360 $X2=0.6210 $Y2=0.0360
r52 31 51 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0360 $X2=0.6750 $Y2=0.0540
r53 2 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6750 $Y=0.1350
+ $X2=0.6750 $Y2=0.1330
r54 14 2 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6750
+ $Y=0.1350 $X2=0.6750 $Y2=0.1350
r55 50 51 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0680 $X2=0.6750 $Y2=0.0540
r56 49 50 1.63233 $w=1.3e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0750 $X2=0.6750 $Y2=0.0680
r57 48 49 0.932759 $w=1.3e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0790 $X2=0.6750 $Y2=0.0750
r58 47 48 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0880 $X2=0.6750 $Y2=0.0790
r59 26 32 1.33376 $w=1.70476e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6750 $Y=0.0970 $X2=0.6750 $Y2=0.1075
r60 26 47 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0970 $X2=0.6750 $Y2=0.0880
r61 44 45 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1205 $X2=0.6750 $Y2=0.1330
r62 43 44 0.867186 $w=1.3625e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.6750 $Y=0.1165 $X2=0.6750 $Y2=0.1205
r63 32 43 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1075 $X2=0.6750 $Y2=0.1165
r64 42 43 6.81353 $w=1.30847e-08 $l=3.89391e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7130 $Y=0.1080 $X2=0.6750 $Y2=0.1165
r65 41 42 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.7445
+ $Y=0.1080 $X2=0.7130 $Y2=0.1080
r66 40 41 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.1080 $X2=0.7445 $Y2=0.1080
r67 27 38 8.26388 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7965 $Y=0.1080 $X2=0.8370 $Y2=0.1080
r68 27 40 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.7965
+ $Y=0.1080 $X2=0.7560 $Y2=0.1080
r69 33 37 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1205 $X2=0.8370 $Y2=0.1330
r70 33 38 1.73456 $w=1.66e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8370 $Y=0.1205 $X2=0.8370 $Y2=0.1080
r71 15 3 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.8370
+ $Y=0.1350 $X2=0.8370 $Y2=0.1350
r72 3 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8370 $Y=0.1350
+ $X2=0.8370 $Y2=0.1330
.ends

.subckt PM_ICGx3_ASAP7_75t_R%NET14 VSS 9 41 42 44 11 13 4 3 12 10 1 14
c1 1 VSS 0.00374789f
c2 3 VSS 0.00716948f
c3 4 VSS 0.0090279f
c4 9 VSS 0.0801723f
c5 10 VSS 0.00631945f
c6 11 VSS 0.00498261f
c7 12 VSS 0.0168337f
c8 13 VSS 0.0107251f
c9 14 VSS 0.00671233f
c10 15 VSS 0.00312913f
c11 16 VSS 0.00353908f
r1 44 43 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r2 11 43 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r3 42 40 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0540 $X2=0.1225 $Y2=0.0540
r4 4 40 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0540 $X2=0.1225 $Y2=0.0540
r5 10 4 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0540 $X2=0.1080 $Y2=0.0540
r6 41 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0540 $X2=0.0935 $Y2=0.0540
r7 3 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0540 $Y2=0.2330
r8 4 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0540
+ $X2=0.1080 $Y2=0.0360
r9 37 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2330 $X2=0.0675 $Y2=0.2330
r10 35 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.2330 $X2=0.0675 $Y2=0.2330
r11 34 35 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2330 $X2=0.0810 $Y2=0.2330
r12 33 34 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2330 $X2=0.1080 $Y2=0.2330
r13 12 16 5.06479 $w=1.46038e-08 $l=2.70046e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1620 $Y=0.2330 $X2=0.1890 $Y2=0.2325
r14 12 33 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2330 $X2=0.1350 $Y2=0.2330
r15 30 31 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.1215 $Y2=0.0360
r16 28 31 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1215 $Y2=0.0360
r17 13 15 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1620 $Y=0.0360 $X2=0.1890 $Y2=0.0360
r18 13 28 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r19 16 26 0.983973 $w=1.77222e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2325 $X2=0.1890 $Y2=0.2235
r20 15 21 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1890 $Y2=0.0575
r21 25 26 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2110 $X2=0.1890 $Y2=0.2235
r22 24 25 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1985 $X2=0.1890 $Y2=0.2110
r23 23 24 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1910 $X2=0.1890 $Y2=0.1985
r24 22 23 9.211 $w=1.3e-08 $l=3.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1515 $X2=0.1890 $Y2=0.1910
r25 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0710 $X2=0.1890 $Y2=0.0575
r26 19 20 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0810 $X2=0.1890 $Y2=0.0710
r27 14 19 5.47996 $w=1.3e-08 $l=2.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1045 $X2=0.1890 $Y2=0.0810
r28 14 22 10.9599 $w=1.3e-08 $l=4.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1045 $X2=0.1890 $Y2=0.1515
r29 9 1 6.2219 $w=1.2115e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1340
r30 1 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1340
+ $X2=0.1890 $Y2=0.1515
r31 3 11 1e-05
.ends

.subckt PM_ICGx3_ASAP7_75t_R%GCLKN VSS 12 13 14 58 59 67 68 71 72 15 17 5 16 3
+ 18 4 19 22 1 21 24 23
c1 1 VSS 0.0142024f
c2 3 VSS 0.00971811f
c3 4 VSS 0.00647354f
c4 5 VSS 0.00935757f
c5 12 VSS 0.0812775f
c6 13 VSS 0.0808804f
c7 14 VSS 0.0807039f
c8 15 VSS 0.00484049f
c9 16 VSS 0.00583673f
c10 17 VSS 0.00581766f
c11 18 VSS 0.013003f
c12 19 VSS 0.00655396f
c13 20 VSS 0.00205696f
c14 21 VSS 0.00291731f
c15 22 VSS 0.00436038f
c16 23 VSS 0.00119776f
c17 24 VSS 0.00137745f
r1 72 70 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.2160 $X2=0.7165 $Y2=0.2160
r2 3 70 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7020 $Y=0.2160 $X2=0.7165 $Y2=0.2160
r3 16 3 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.2160 $X2=0.7020 $Y2=0.2160
r4 71 16 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.2160 $X2=0.6875 $Y2=0.2160
r5 68 66 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8270 $Y=0.2160 $X2=0.8245 $Y2=0.2160
r6 5 66 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8100 $Y=0.2160 $X2=0.8245 $Y2=0.2160
r7 17 5 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.2160 $X2=0.8100 $Y2=0.2160
r8 67 17 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.2160 $X2=0.7955 $Y2=0.2160
r9 3 63 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7020 $Y=0.2160
+ $X2=0.7020 $Y2=0.2310
r10 5 60 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8100 $Y=0.2160
+ $X2=0.8100 $Y2=0.2310
r11 63 64 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.2310 $X2=0.7380 $Y2=0.2310
r12 60 61 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.2310 $X2=0.8235 $Y2=0.2310
r13 18 60 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.2310 $X2=0.8100 $Y2=0.2310
r14 18 64 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.2310 $X2=0.7380 $Y2=0.2310
r15 58 57 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.0675 $X2=0.7705 $Y2=0.0675
r16 4 57 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7560 $Y=0.0675 $X2=0.7705 $Y2=0.0675
r17 15 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7415 $Y=0.0675 $X2=0.7560 $Y2=0.0675
r18 59 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.0675 $X2=0.7415 $Y2=0.0675
r19 54 61 1.20242 $w=1.425e-08 $l=1.54434e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8370 $Y=0.2235 $X2=0.8235 $Y2=0.2310
r20 53 54 2.01858 $w=1.37895e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.8370 $Y=0.2140 $X2=0.8370 $Y2=0.2235
r21 52 53 2.37574 $w=1.49231e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8370 $Y=0.2010 $X2=0.8370 $Y2=0.2140
r22 22 52 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1920 $X2=0.8370 $Y2=0.2010
r23 4 50 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7560 $Y=0.0675
+ $X2=0.7560 $Y2=0.0720
r24 20 24 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8640 $Y=0.1970 $X2=0.8910 $Y2=0.1970
r25 20 22 4.60559 $w=1.39091e-08 $l=2.74591e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8640 $Y=0.1970 $X2=0.8370 $Y2=0.1920
r26 50 51 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.0720 $X2=0.7965 $Y2=0.0720
r27 48 51 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.0720 $X2=0.7965 $Y2=0.0720
r28 47 48 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.8625
+ $Y=0.0720 $X2=0.8370 $Y2=0.0720
r29 19 23 0.79938 $w=1.72857e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8805 $Y=0.0720 $X2=0.8910 $Y2=0.0720
r30 19 47 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8805
+ $Y=0.0720 $X2=0.8625 $Y2=0.0720
r31 24 44 5.22999 $w=1.59898e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8910 $Y=0.1970 $X2=0.8910 $Y2=0.1675
r32 23 43 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.0720 $X2=0.8910 $Y2=0.0900
r33 14 39 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=0.9990
+ $Y=0.1350 $X2=0.9990 $Y2=0.1360
r34 13 33 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=0.9450
+ $Y=0.1350 $X2=0.9450 $Y2=0.1360
r35 42 44 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1460 $X2=0.8910 $Y2=0.1675
r36 41 42 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1360 $X2=0.8910 $Y2=0.1460
r37 21 41 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1130 $X2=0.8910 $Y2=0.1360
r38 21 43 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1130 $X2=0.8910 $Y2=0.0900
r39 37 39 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9865 $Y=0.1360 $X2=0.9990 $Y2=0.1360
r40 36 37 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9720 $Y=0.1360 $X2=0.9865 $Y2=0.1360
r41 34 36 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9575 $Y=0.1360 $X2=0.9720 $Y2=0.1360
r42 33 34 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9450 $Y=0.1360 $X2=0.9575 $Y2=0.1360
r43 31 33 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9325 $Y=0.1360 $X2=0.9450 $Y2=0.1360
r44 30 31 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9180 $Y=0.1360 $X2=0.9325 $Y2=0.1360
r45 29 30 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9035 $Y=0.1360 $X2=0.9180 $Y2=0.1360
r46 27 29 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.9005 $Y=0.1360 $X2=0.9035 $Y2=0.1360
r47 26 27 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.8910
+ $Y=0.1360 $X2=0.9005 $Y2=0.1360
r48 26 41 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8910 $Y=0.1360
+ $X2=0.8910 $Y2=0.1360
r49 1 26 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.8815
+ $Y=0.1360 $X2=0.8910 $Y2=0.1360
r50 1 28 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.8815
+ $Y=0.1360 $X2=0.8805 $Y2=0.1360
r51 12 26 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.8910 $Y=0.1350 $X2=0.8910 $Y2=0.1360
r52 12 28 0.610027 $w=2.16919e-07 $l=1.05475e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.8910 $Y=0.1350 $X2=0.8805 $Y2=0.1360
r53 12 29 1.79147 $w=1.8466e-07 $l=1.25399e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.8910 $Y=0.1350 $X2=0.9035 $Y2=0.1360
.ends

.subckt PM_ICGx3_ASAP7_75t_R%CLKN VSS 9 53 55 10 13 18 3 15 12 1 11 17 14 16 4
c1 1 VSS 9.81683e-20
c2 3 VSS 0.00618855f
c3 4 VSS 0.00786156f
c4 9 VSS 0.00447213f
c5 10 VSS 0.00617799f
c6 11 VSS 0.00620482f
c7 12 VSS 0.000529362f
c8 13 VSS 0.00120981f
c9 14 VSS 0.00264871f
c10 15 VSS 0.000644133f
c11 16 VSS 0.00085415f
c12 17 VSS 0.00632271f
c13 18 VSS 0.00872721f
r1 55 54 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.2025 $X2=0.6085 $Y2=0.2025
r2 11 54 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5960 $Y=0.2025 $X2=0.6085 $Y2=0.2025
r3 53 52 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.0675 $X2=0.6085 $Y2=0.0675
r4 10 52 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5960 $Y=0.0675 $X2=0.6085 $Y2=0.0675
r5 4 46 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2295
+ $X2=0.5940 $Y2=0.2320
r6 3 43 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0605
+ $X2=0.5940 $Y2=0.0860
r7 45 46 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5810
+ $Y=0.2320 $X2=0.5940 $Y2=0.2320
r8 17 41 1.03499 $w=1.77368e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.5680 $Y=0.2320 $X2=0.5680 $Y2=0.2225
r9 17 45 1.85116 $w=1.64615e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5680 $Y=0.2320 $X2=0.5810 $Y2=0.2320
r10 42 43 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5810
+ $Y=0.0860 $X2=0.5940 $Y2=0.0860
r11 16 38 3.36689 $w=1.53077e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5680 $Y=0.0860 $X2=0.5680 $Y2=0.1055
r12 16 42 1.85116 $w=1.64615e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5680 $Y=0.0860 $X2=0.5810 $Y2=0.0860
r13 40 41 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5680
+ $Y=0.2100 $X2=0.5680 $Y2=0.2225
r14 39 40 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5680
+ $Y=0.1970 $X2=0.5680 $Y2=0.2100
r15 37 39 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5680
+ $Y=0.1880 $X2=0.5680 $Y2=0.1970
r16 13 37 9.32759 $w=1.3e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.5680
+ $Y=0.1480 $X2=0.5680 $Y2=0.1880
r17 13 38 9.91056 $w=1.3e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5680
+ $Y=0.1480 $X2=0.5680 $Y2=0.1055
r18 35 37 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.5680 $Y=0.1890
+ $X2=0.5680 $Y2=0.1880
r19 34 35 30.0815 $w=1.3e-08 $l=1.29e-07 $layer=M2 $thickness=3.6e-08 $X=0.4390
+ $Y=0.1890 $X2=0.5680 $Y2=0.1890
r20 33 34 30.0815 $w=1.3e-08 $l=1.29e-07 $layer=M2 $thickness=3.6e-08 $X=0.3100
+ $Y=0.1890 $X2=0.4390 $Y2=0.1890
r21 18 33 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.2985
+ $Y=0.1890 $X2=0.3100 $Y2=0.1890
r22 31 33 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.3145 $Y=0.1890
+ $X2=0.3100 $Y2=0.1890
r23 30 31 1.51573 $w=1.3e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3080
+ $Y=0.1890 $X2=0.3145 $Y2=0.1890
r24 29 30 0.721491 $w=1.57778e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.3035 $Y=0.1890 $X2=0.3080 $Y2=0.1890
r25 15 29 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2945
+ $Y=0.1890 $X2=0.3035 $Y2=0.1890
r26 27 29 4.68572 $w=1.35814e-08 $l=2.87446e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1610 $X2=0.3035 $Y2=0.1890
r27 26 27 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1330 $X2=0.2970 $Y2=0.1610
r28 25 26 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1215 $X2=0.2970 $Y2=0.1330
r29 12 25 3.96423 $w=1.3e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1045 $X2=0.2970 $Y2=0.1215
r30 12 14 4.29965 $w=1.49149e-08 $l=2.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1045 $X2=0.2970 $Y2=0.0810
r31 1 22 2.88023 $w=2.1e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.2970
+ $Y=0.1335 $X2=0.2970 $Y2=0.1335
r32 1 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1335
+ $X2=0.2970 $Y2=0.1330
r33 9 22 0.314665 $w=2.27e-07 $l=1.5e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2970 $Y2=0.1335
r34 4 11 1e-05
r35 3 10 1e-05
.ends

.subckt PM_ICGx3_ASAP7_75t_R%CLK VSS 49 10 11 12 13 14 23 1 15 21 20 16 8 17 3
+ 2 19 22 4 18
c1 1 VSS 0.00383292f
c2 2 VSS 0.00186666f
c3 3 VSS 0.00738049f
c4 4 VSS 0.00893638f
c5 8 VSS 0.00400423f
c6 10 VSS 0.00632478f
c7 11 VSS 0.0062577f
c8 12 VSS 0.0820853f
c9 13 VSS 0.0342495f
c10 14 VSS 0.0342998f
c11 15 VSS 0.00473339f
c12 16 VSS 0.00463287f
c13 17 VSS 0.00488878f
c14 18 VSS 0.00226697f
c15 19 VSS 0.00195735f
c16 20 VSS 0.00386868f
c17 21 VSS 0.00246759f
c18 22 VSS 0.00242725f
c19 23 VSS 0.00603415f
r1 2 78 3.16825 $w=2.1e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.3520
+ $Y=0.1335 $X2=0.3555 $Y2=0.1335
r2 11 2 3.48292 $w=1.19095e-07 $l=1.80278e-09 $layer=LIG $thickness=5.18095e-08
+ $X=0.3510 $Y=0.1350 $X2=0.3520 $Y2=0.1335
r3 77 78 4.91375 $w=2.12e-08 $l=1.5e-09 $layer=LISD $thickness=2.7e-08
+ $X=0.3570 $Y=0.1335 $X2=0.3555 $Y2=0.1335
r4 76 77 11.4654 $w=2.12e-08 $l=2.1e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.3780 $Y=0.1335 $X2=0.3570 $Y2=0.1335
r5 75 76 7.37062 $w=2.12e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.3915 $Y=0.1335 $X2=0.3780 $Y2=0.1335
r6 8 73 5.7327 $w=2.12e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08 $X=0.3945
+ $Y=0.1335 $X2=0.4050 $Y2=0.1335
r7 8 75 1.63792 $w=2.12e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.3945
+ $Y=0.1335 $X2=0.3915 $Y2=0.1335
r8 1 62 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1335
+ $X2=0.2430 $Y2=0.1330
r9 10 1 3.19489 $w=1.24e-07 $l=1.5e-09 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1335
r10 69 70 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1340 $X2=0.4050 $Y2=0.1435
r11 69 73 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4050 $Y=0.1340
+ $X2=0.4050 $Y2=0.1335
r12 19 20 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1530 $X2=0.4230 $Y2=0.1530
r13 19 70 1.03499 $w=1.77368e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.1530 $X2=0.4050 $Y2=0.1435
r14 63 64 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1430 $X2=0.2430 $Y2=0.1530
r15 62 63 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1330 $X2=0.2430 $Y2=0.1430
r16 15 62 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1215 $X2=0.2430 $Y2=0.1330
r17 20 54 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4230 $Y=0.1530
+ $X2=0.4230 $Y2=0.1530
r18 3 46 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6210 $Y=0.1350
+ $X2=0.6210 $Y2=0.1330
r19 12 3 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1350
r20 57 58 7.22888 $w=1.3e-08 $l=3.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1530 $X2=0.2740 $Y2=0.1530
r21 57 64 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.2430 $Y=0.1530
+ $X2=0.2430 $Y2=0.1530
r22 54 55 19.5879 $w=1.3e-08 $l=8.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.4230
+ $Y=0.1530 $X2=0.5070 $Y2=0.1530
r23 53 54 15.8569 $w=1.3e-08 $l=6.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.3550
+ $Y=0.1530 $X2=0.4230 $Y2=0.1530
r24 53 58 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.3550
+ $Y=0.1530 $X2=0.2740 $Y2=0.1530
r25 50 51 4.25571 $w=1.3e-08 $l=1.83e-08 $layer=M2 $thickness=3.6e-08 $X=0.6027
+ $Y=0.1530 $X2=0.6210 $Y2=0.1530
r26 49 50 2.2736 $w=1.3e-08 $l=9.7e-09 $layer=M2 $thickness=3.6e-08 $X=0.5930
+ $Y=0.1530 $X2=0.6027 $Y2=0.1530
r27 49 23 1.34084 $w=1.3e-08 $l=5.8e-09 $layer=M2 $thickness=3.6e-08 $X=0.5930
+ $Y=0.1530 $X2=0.5872 $Y2=0.1530
r28 23 55 18.7135 $w=1.3e-08 $l=8.02e-08 $layer=M2 $thickness=3.6e-08 $X=0.5872
+ $Y=0.1530 $X2=0.5070 $Y2=0.1530
r29 47 48 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1430 $X2=0.6210 $Y2=0.1455
r30 46 47 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1330 $X2=0.6210 $Y2=0.1430
r31 16 44 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1545 $X2=0.6210 $Y2=0.1700
r32 16 48 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1545 $X2=0.6210 $Y2=0.1455
r33 16 51 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.6210 $Y=0.1545
+ $X2=0.6210 $Y2=0.1530
r34 21 43 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.1870 $X2=0.6480 $Y2=0.1870
r35 21 44 2.31511 $w=1.81882e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.1870 $X2=0.6210 $Y2=0.1700
r36 42 43 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1870 $X2=0.6480 $Y2=0.1870
r37 41 42 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6860
+ $Y=0.1870 $X2=0.6750 $Y2=0.1870
r38 17 22 7.38932 $w=1.37246e-08 $l=3.87072e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7175 $Y=0.1870 $X2=0.7560 $Y2=0.1830
r39 17 41 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.7175
+ $Y=0.1870 $X2=0.6860 $Y2=0.1870
r40 22 38 1.32639 $w=1.59412e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.7560 $Y=0.1830 $X2=0.7560 $Y2=0.1745
r41 13 33 2.92627 $w=1.245e-07 $l=2.7e-08 $layer=LIG $thickness=5.2e-08
+ $X=0.7290 $Y=0.1350 $X2=0.7290 $Y2=0.1620
r42 37 38 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.1620 $X2=0.7560 $Y2=0.1745
r43 36 37 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.1500 $X2=0.7560 $Y2=0.1620
r44 18 36 1.28254 $w=1.3e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.1445 $X2=0.7560 $Y2=0.1500
r45 31 33 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7415 $Y=0.1620 $X2=0.7290 $Y2=0.1620
r46 30 31 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7560 $Y=0.1620 $X2=0.7415 $Y2=0.1620
r47 30 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7560 $Y=0.1620
+ $X2=0.7560 $Y2=0.1620
r48 29 30 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7705 $Y=0.1620 $X2=0.7560 $Y2=0.1620
r49 4 28 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.7830
+ $Y=0.1620 $X2=0.7830 $Y2=0.1620
r50 4 29 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7830 $Y=0.1620 $X2=0.7705 $Y2=0.1620
r51 4 35 2.90696 $w=2.1681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7830 $Y=0.1620 $X2=0.7935 $Y2=0.1620
r52 28 29 1.47681 $w=1.53e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7830 $Y=0.1620 $X2=0.7705 $Y2=0.1620
r53 28 35 0.295362 $w=1.53e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7830 $Y=0.1620 $X2=0.7935 $Y2=0.1620
r54 14 28 0.314665 $w=2.27e-07 $l=2.7e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.7830 $Y=0.1350 $X2=0.7830 $Y2=0.1620
.ends


*
.SUBCKT ICGx3_ASAP7_75t_R VSS VDD ENA SE CLK GCLK
*
* VSS VSS
* VDD VDD
* ENA ENA
* SE SE
* CLK CLK
* GCLK GCLK
*
*

MM19 N_MM19_d N_MM19_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM27 N_MM27_d N_MM18_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM10_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM6 N_MM6_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM20 N_MM20_d N_MM21_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM14 N_MM14_d N_MM0_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM16_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM13 N_MM13_d N_MM13_g N_MM13_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM12 N_MM12_d N_MM12_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24 N_MM24_d N_MM24_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@3 N_MM24@3_d N_MM24@3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@2 N_MM24@2_d N_MM24@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM26 N_MM26_d N_MM19_g N_MM26_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM18 N_MM18_d N_MM18_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM21 N_MM21_d N_MM21_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM16 N_MM16_d N_MM16_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM16@2 N_MM16@2_d N_MM13_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM0@2 N_MM0@2_d N_MM12_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM25 N_MM25_d N_MM24_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@3 N_MM25@3_d N_MM24@3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@2 N_MM25@2_d N_MM24@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "ICGx3_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "ICGx3_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_ICGx3_ASAP7_75t_R%NOS1 VSS N_MM26_s N_MM18_d N_NOS1_1
+ PM_ICGx3_ASAP7_75t_R%NOS1
cc_1 N_NOS1_1 N_MM19_g 0.0125258f
cc_2 N_NOS1_1 N_MM18_g 0.0125785f
x_PM_ICGx3_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_ICGx3_ASAP7_75t_R%noxref_19
cc_3 N_noxref_19_1 N_MM19_g 0.00394297f
cc_4 N_noxref_19_1 N_NET14_10 0.00040021f
x_PM_ICGx3_ASAP7_75t_R%ENA VSS ENA N_MM19_g N_ENA_1 N_ENA_4
+ PM_ICGx3_ASAP7_75t_R%ENA
x_PM_ICGx3_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_ICGx3_ASAP7_75t_R%noxref_20
cc_5 N_noxref_20_1 N_MM19_g 0.00393678f
cc_6 N_noxref_20_1 N_NET14_11 0.0276623f
cc_7 N_noxref_20_1 N_noxref_19_1 0.00208841f
x_PM_ICGx3_ASAP7_75t_R%SE VSS SE N_MM18_g N_SE_1 N_SE_4 PM_ICGx3_ASAP7_75t_R%SE
cc_8 N_SE_1 N_ENA_1 0.00169567f
cc_9 N_SE_4 N_ENA_4 0.00508575f
cc_10 N_MM18_g N_MM19_g 0.00985319f
x_PM_ICGx3_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_ICGx3_ASAP7_75t_R%noxref_25
cc_11 N_noxref_25_1 N_MM24@2_g 0.00145528f
cc_12 N_noxref_25_1 N_GCLK_14 0.0378538f
x_PM_ICGx3_ASAP7_75t_R%noxref_26 VSS N_noxref_26_1
+ PM_ICGx3_ASAP7_75t_R%noxref_26
cc_13 N_noxref_26_1 N_MM24@2_g 0.00146208f
cc_14 N_noxref_26_1 N_GCLK_16 0.0376114f
cc_15 N_noxref_26_1 N_noxref_25_1 0.00177022f
x_PM_ICGx3_ASAP7_75t_R%GCLK VSS GCLK N_MM24_d N_MM24@3_d N_MM24@2_d N_MM25_d
+ N_MM25@3_d N_MM25@2_d N_GCLK_13 N_GCLK_17 N_GCLK_3 N_GCLK_15 N_GCLK_4
+ N_GCLK_1 N_GCLK_2 N_GCLK_18 N_GCLK_16 N_GCLK_14 PM_ICGx3_ASAP7_75t_R%GCLK
cc_16 N_GCLK_13 N_GCLKN_1 0.00113355f
cc_17 N_GCLK_13 N_MM24@2_g 0.0008843f
cc_18 N_GCLK_17 N_GCLKN_19 0.000835707f
cc_19 N_GCLK_3 N_MM24@2_g 0.00087479f
cc_20 N_GCLK_15 N_MM24@3_g 0.0309364f
cc_21 N_GCLK_4 N_MM24@2_g 0.000898769f
cc_22 N_GCLK_1 N_GCLKN_21 0.00164441f
cc_23 N_GCLK_1 N_MM24@3_g 0.00224994f
cc_24 N_GCLK_2 N_MM24@3_g 0.00238104f
cc_25 N_GCLK_18 N_GCLKN_24 0.0025512f
cc_26 N_GCLK_17 N_GCLKN_23 0.00327584f
cc_27 N_GCLK_16 N_MM24@2_g 0.0148656f
cc_28 N_GCLK_15 N_GCLKN_1 0.00673152f
cc_29 N_GCLK_14 N_MM24@2_g 0.0527291f
cc_30 N_GCLK_13 N_MM24_g 0.0371335f
cc_31 N_GCLK_13 N_MM24@3_g 0.0692619f
x_PM_ICGx3_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_ICGx3_ASAP7_75t_R%noxref_22
cc_32 N_noxref_22_1 N_CLKN_11 0.000956656f
cc_33 N_noxref_22_1 N_MS_11 0.0170564f
cc_34 N_noxref_22_1 N_MM7_g 0.00577904f
cc_35 N_noxref_22_1 N_noxref_21_1 0.00153657f
x_PM_ICGx3_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_ICGx3_ASAP7_75t_R%noxref_21
cc_36 N_noxref_21_1 N_CLKN_10 0.000837518f
cc_37 N_noxref_21_1 N_MS_3 0.00100914f
cc_38 N_noxref_21_1 N_MS_10 0.0169534f
cc_39 N_noxref_21_1 N_MM7_g 0.00534655f
x_PM_ICGx3_ASAP7_75t_R%NET056 VSS N_MM14_d N_MM2_s N_NET056_1
+ PM_ICGx3_ASAP7_75t_R%NET056
cc_40 N_NET056_1 N_MM16_g 0.0174349f
cc_41 N_NET056_1 N_MM0_g 0.0172741f
x_PM_ICGx3_ASAP7_75t_R%PD3 VSS N_MM9_s N_MM8_d N_PD3_3 N_PD3_1
+ PM_ICGx3_ASAP7_75t_R%PD3
cc_42 N_PD3_3 N_MM9_g 0.0146784f
cc_43 N_PD3_3 N_MM11_g 0.0162408f
cc_44 N_PD3_1 N_MH_22 0.000207302f
cc_45 N_PD3_1 N_MH_16 0.000611638f
cc_46 N_PD3_1 N_MH_24 0.000293363f
cc_47 N_PD3_1 N_MH_8 0.00212236f
x_PM_ICGx3_ASAP7_75t_R%PU1 VSS N_MM3_d N_MM1_s N_PU1_3 N_PU1_1
+ PM_ICGx3_ASAP7_75t_R%PU1
cc_48 N_PU1_3 N_NET14_1 0.000627842f
cc_49 N_PU1_3 N_MM3_g 0.0349004f
cc_50 N_PU1_3 N_CLK_15 0.000334715f
cc_51 N_PU1_3 N_CLK_1 0.000513648f
cc_52 N_PU1_3 N_MM1_g 0.0336029f
cc_53 N_PU1_1 N_MH_18 0.00109778f
cc_54 N_PU1_1 N_MH_7 0.00288975f
x_PM_ICGx3_ASAP7_75t_R%MS VSS N_MM11_g N_MM6_d N_MM7_d N_MS_1 N_MS_12 N_MS_13
+ N_MS_15 N_MS_3 N_MS_14 N_MS_4 N_MS_11 N_MS_10 PM_ICGx3_ASAP7_75t_R%MS
cc_55 N_MM11_g N_CLK_20 0.000217535f
cc_56 N_MM11_g N_CLK_23 0.000125382f
cc_57 N_MM11_g N_CLK_8 0.00294031f
cc_58 N_MS_1 N_CLK_19 0.000552116f
cc_59 N_MS_1 N_CLK_8 0.00153715f
cc_60 N_MS_12 N_CLK_20 0.000626225f
cc_61 N_MS_13 N_CLK_23 0.00150955f
cc_62 N_MS_12 N_CLK_23 0.001564f
cc_63 N_MS_12 N_CLK_19 0.00255782f
cc_64 N_MM11_g N_MM9_g 0.0131996f
cc_65 N_MS_13 N_CLKN_11 0.000122571f
cc_66 N_MS_13 N_CLKN_16 0.000223033f
cc_67 N_MS_15 N_CLKN_3 0.00024744f
cc_68 N_MS_3 N_CLKN_16 0.000253119f
cc_69 N_MS_13 N_CLKN_4 0.000275436f
cc_70 N_MS_14 N_CLKN_17 0.000855618f
cc_71 N_MS_15 N_CLKN_16 0.000951897f
cc_72 N_MS_14 N_CLKN_18 0.00148628f
cc_73 N_MS_13 N_CLKN_13 0.00669115f
x_PM_ICGx3_ASAP7_75t_R%PD1 VSS N_MM5_d N_MM4_s N_PD1_4 N_PD1_5 N_PD1_1
+ PM_ICGx3_ASAP7_75t_R%PD1
cc_74 N_PD1_4 N_NET14_1 0.000768641f
cc_75 N_PD1_4 N_MM3_g 0.0359403f
cc_76 N_PD1_5 N_CLK_1 0.00231353f
cc_77 N_PD1_5 N_MM1_g 0.0731939f
cc_78 N_PD1_5 N_CLKN_1 0.000683141f
cc_79 N_PD1_5 N_CLKN_14 0.00273042f
cc_80 N_PD1_5 N_MM10_g 0.0334545f
cc_81 N_PD1_1 N_MH_8 0.00133102f
cc_82 N_PD1_1 N_MH_16 0.00293317f
x_PM_ICGx3_ASAP7_75t_R%NET059 VSS N_MM13_s N_MM12_d N_NET059_1
+ PM_ICGx3_ASAP7_75t_R%NET059
cc_83 N_NET059_1 N_MM13_g 0.0173246f
cc_84 N_NET059_1 N_MM12_g 0.0173168f
x_PM_ICGx3_ASAP7_75t_R%PD2 VSS N_MM10_s N_MM11_d N_PD2_5 N_PD2_4 N_PD2_1
+ PM_ICGx3_ASAP7_75t_R%PD2
cc_85 N_PD2_5 N_CLK_8 0.000220944f
cc_86 N_PD2_4 N_MM9_g 0.00732296f
cc_87 N_PD2_1 N_MM9_g 0.0009939f
cc_88 N_PD2_5 N_MM9_g 0.0237233f
cc_89 N_PD2_1 N_MM10_g 0.000492671f
cc_90 N_PD2_4 N_MM10_g 0.0149714f
cc_91 N_PD2_5 N_MM11_g 0.0149321f
cc_92 N_PD2_1 N_MH_22 9.53537e-20
cc_93 N_PD2_1 N_MH_7 0.000117211f
cc_94 N_PD2_1 N_MH_23 0.000256152f
cc_95 N_PD2_1 N_MH_25 0.000296431f
cc_96 N_PD2_4 N_MH_18 0.000643006f
cc_97 N_PD2_1 N_MH_20 0.000491765f
cc_98 N_PD2_4 N_MH_7 0.000618537f
cc_99 N_PD2_1 N_MH_30 0.002704f
x_PM_ICGx3_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_ICGx3_ASAP7_75t_R%noxref_24
cc_100 N_noxref_24_1 N_MM21_g 0.00136834f
cc_101 N_noxref_24_1 N_CLKN_4 0.00041051f
cc_102 N_noxref_24_1 N_CLKN_11 0.0373735f
cc_103 N_noxref_24_1 N_MS_11 0.00053837f
cc_104 N_noxref_24_1 N_noxref_21_1 0.000473227f
cc_105 N_noxref_24_1 N_noxref_22_1 0.00777077f
cc_106 N_noxref_24_1 N_noxref_23_1 0.00123137f
x_PM_ICGx3_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_ICGx3_ASAP7_75t_R%noxref_23
cc_107 N_noxref_23_1 N_MM21_g 0.00136327f
cc_108 N_noxref_23_1 N_CLKN_10 0.0376459f
cc_109 N_noxref_23_1 N_MS_10 0.000573044f
cc_110 N_noxref_23_1 N_noxref_21_1 0.00773065f
cc_111 N_noxref_23_1 N_noxref_22_1 0.000477267f
x_PM_ICGx3_ASAP7_75t_R%MH VSS N_MM7_g N_MM0_g N_MM12_g N_MM4_d N_MM9_d N_MM1_d
+ N_MM10_d N_MH_23 N_MH_7 N_MH_21 N_MH_29 N_MH_19 N_MH_17 N_MH_27 N_MH_32
+ N_MH_33 N_MH_18 N_MH_3 N_MH_1 N_MH_25 N_MH_26 N_MH_20 N_MH_22 N_MH_24 N_MH_16
+ N_MH_8 N_MH_2 N_MH_30 N_MH_31 PM_ICGx3_ASAP7_75t_R%MH
cc_112 N_MH_23 N_CLK_19 7.89505e-20
cc_113 N_MH_7 N_CLK_15 0.000840224f
cc_114 N_MH_21 N_MM9_g 0.000133524f
cc_115 N_MH_29 N_CLK_19 0.000143071f
cc_116 N_MH_19 N_MM1_g 0.00014953f
cc_117 N_MH_17 N_MM9_g 0.000175721f
cc_118 N_MH_27 N_CLK_22 0.000201848f
cc_119 N_MH_7 N_CLK_1 0.000204324f
cc_120 N_MH_32 N_CLK_16 0.00305632f
cc_121 N_MH_33 N_CLK_4 0.000243122f
cc_122 N_MH_18 N_MM1_g 0.0338941f
cc_123 N_MH_3 N_CLK_4 0.000266968f
cc_124 N_MH_1 N_CLK_8 0.000271258f
cc_125 N_MH_1 N_CLK_20 0.000305803f
cc_126 N_MH_25 N_CLK_20 0.00476149f
cc_127 N_MH_26 N_CLK_16 0.000363298f
cc_128 N_MH_27 N_CLK_4 0.000401496f
cc_129 N_MH_20 N_CLK_15 0.000487313f
cc_130 N_MH_22 N_CLK_8 0.00250082f
cc_131 N_MM7_g N_CLK_8 0.00054433f
cc_132 N_MH_3 N_MM13_g 0.000546272f
cc_133 N_MH_18 N_CLK_1 0.000569951f
cc_134 N_MH_24 N_CLK_23 0.000690775f
cc_135 N_MH_16 N_CLK_2 0.000886988f
cc_136 N_MH_8 N_MM9_g 0.00101642f
cc_137 N_MH_7 N_MM1_g 0.0011796f
cc_138 N_MH_2 N_CLK_3 0.00305765f
cc_139 N_MH_25 N_CLK_19 0.00140162f
cc_140 N_MH_32 N_CLK_17 0.0015053f
cc_141 N_MM12_g N_CLK_4 0.00166613f
cc_142 N_MM0_g N_MM21_g 0.00166641f
cc_143 N_MH_25 N_CLK_23 0.00230474f
cc_144 N_MH_27 N_CLK_18 0.00377593f
cc_145 N_MH_22 N_CLK_19 0.00383142f
cc_146 N_MM12_g N_MM13_g 0.00715355f
cc_147 N_MM0_g N_MM16_g 0.00886723f
cc_148 N_MH_16 N_MM9_g 0.0366474f
cc_149 N_MM0_g N_MM10_g 0.000126632f
cc_150 N_MH_27 N_MM10_g 8.92992e-20
cc_151 N_MM7_g N_MM10_g 9.38751e-20
cc_152 N_MH_17 N_MM10_g 0.000144983f
cc_153 N_MH_32 N_CLKN_16 0.000150038f
cc_154 N_MH_19 N_MM10_g 0.000166264f
cc_155 N_MH_8 N_CLKN_14 0.000186868f
cc_156 N_MH_7 N_CLKN_15 0.000193659f
cc_157 N_MH_30 N_CLKN_15 0.000197599f
cc_158 N_MH_26 N_CLKN_16 0.00021494f
cc_159 N_MH_25 N_CLKN_13 0.000249005f
cc_160 N_MH_24 N_CLKN_3 0.00111962f
cc_161 N_MH_18 N_MM10_g 0.0166804f
cc_162 N_MH_20 N_CLKN_15 0.00477986f
cc_163 N_MH_23 N_CLKN_15 0.000541385f
cc_164 N_MH_29 N_CLKN_15 0.000688789f
cc_165 N_MH_8 N_CLKN_1 0.000701545f
cc_166 N_MH_8 N_MM10_g 0.00133706f
cc_167 N_MH_7 N_MM10_g 0.00142321f
cc_168 N_MH_16 N_CLKN_1 0.00148257f
cc_169 N_MH_21 N_CLKN_14 0.0019042f
cc_170 N_MH_25 N_CLKN_18 0.00329351f
cc_171 N_MH_22 N_CLKN_12 0.00379305f
cc_172 N_MH_24 N_CLKN_16 0.0043582f
cc_173 N_MH_16 N_MM10_g 0.0536179f
cc_174 N_MH_8 N_MM11_g 0.000202446f
cc_175 N_MH_24 N_MM11_g 0.000315363f
cc_176 N_MH_1 N_MS_4 0.00197807f
cc_177 N_MM7_g N_MS_1 0.000552093f
cc_178 N_MH_24 N_MS_1 0.000727436f
cc_179 N_MH_1 N_MS_11 0.0012631f
cc_180 N_MH_22 N_MS_12 0.00130815f
cc_181 N_MH_25 N_MS_13 0.0013873f
cc_182 N_MM7_g N_MS_3 0.00170061f
cc_183 N_MH_25 N_MS_14 0.00239907f
cc_184 N_MM7_g N_MS_10 0.00643105f
cc_185 N_MM7_g N_MS_11 0.00675895f
cc_186 N_MH_24 N_MS_12 0.00369066f
cc_187 N_MH_24 N_MS_15 0.005497f
cc_188 N_MM7_g N_MM11_g 0.0297137f
x_PM_ICGx3_ASAP7_75t_R%NET14 VSS N_MM3_g N_MM19_d N_MM27_d N_MM26_d N_NET14_11
+ N_NET14_13 N_NET14_4 N_NET14_3 N_NET14_12 N_NET14_10 N_NET14_1 N_NET14_14
+ PM_ICGx3_ASAP7_75t_R%NET14
cc_189 N_NET14_11 N_ENA_1 0.000579346f
cc_190 N_NET14_13 N_ENA_4 0.000723213f
cc_191 N_NET14_4 N_MM19_g 0.000750777f
cc_192 N_NET14_3 N_MM19_g 0.00108943f
cc_193 N_NET14_12 N_ENA_4 0.00143518f
cc_194 N_NET14_4 N_ENA_4 0.00303545f
cc_195 N_NET14_11 N_MM19_g 0.0111053f
cc_196 N_NET14_10 N_MM19_g 0.0403051f
cc_197 N_NET14_1 N_MM18_g 0.00097167f
cc_198 N_NET14_13 N_SE_4 0.00103662f
cc_199 N_NET14_1 N_SE_1 0.00119135f
cc_200 N_NET14_12 N_SE_4 0.00121381f
cc_201 N_NET14_10 N_MM18_g 0.0109236f
cc_202 N_NET14_14 N_SE_4 0.00753965f
cc_203 N_MM3_g N_MM18_g 0.0186725f
x_PM_ICGx3_ASAP7_75t_R%GCLKN VSS N_MM24_g N_MM24@3_g N_MM24@2_g N_MM13_d
+ N_MM2_d N_MM16@2_d N_MM0@2_d N_MM0_d N_MM16_d N_GCLKN_15 N_GCLKN_17 N_GCLKN_5
+ N_GCLKN_16 N_GCLKN_3 N_GCLKN_18 N_GCLKN_4 N_GCLKN_19 N_GCLKN_22 N_GCLKN_1
+ N_GCLKN_21 N_GCLKN_24 N_GCLKN_23 PM_ICGx3_ASAP7_75t_R%GCLKN
cc_204 N_GCLKN_15 N_CLK_4 9.42065e-20
cc_205 N_GCLKN_15 N_CLK_22 0.000418687f
cc_206 N_GCLKN_15 N_CLK_23 0.000176269f
cc_207 N_GCLKN_15 N_CLK_18 0.000285673f
cc_208 N_GCLKN_17 N_MM13_g 0.011333f
cc_209 N_GCLKN_5 N_CLK_4 0.000341215f
cc_210 N_GCLKN_16 N_MM16_g 0.011547f
cc_211 N_GCLKN_3 N_CLK_17 0.000420541f
cc_212 N_GCLKN_18 N_CLK_18 0.000488618f
cc_213 N_GCLKN_5 N_MM13_g 0.000859503f
cc_214 N_GCLKN_3 N_MM16_g 0.00126558f
cc_215 N_GCLKN_4 N_MM13_g 0.00150636f
cc_216 N_GCLKN_17 N_CLK_4 0.00246685f
cc_217 N_GCLKN_18 N_CLK_17 0.00261615f
cc_218 N_GCLKN_18 N_CLK_22 0.00384598f
cc_219 N_GCLKN_15 N_MM16_g 0.0332745f
cc_220 N_GCLKN_15 N_MM13_g 0.0654146f
cc_221 N_GCLKN_16 N_MH_32 0.000115251f
cc_222 N_GCLKN_16 N_MH_2 0.000447009f
cc_223 N_GCLKN_16 N_MH_31 0.000154528f
cc_224 N_GCLKN_16 N_MH_33 0.000496179f
cc_225 N_GCLKN_15 N_MM12_g 0.00030072f
cc_226 N_GCLKN_17 N_MM12_g 0.0112376f
cc_227 N_GCLKN_19 N_MH_26 0.000370132f
cc_228 N_GCLKN_5 N_MM12_g 0.000395902f
cc_229 N_GCLKN_3 N_MM0_g 0.000411282f
cc_230 N_GCLKN_22 N_MH_33 0.00049674f
cc_231 N_GCLKN_4 N_MH_27 0.00182649f
cc_232 N_GCLKN_1 N_MH_3 0.00245999f
cc_233 N_GCLKN_19 N_MH_33 0.00135518f
cc_234 N_GCLKN_21 N_MH_33 0.00270046f
cc_235 N_GCLKN_19 N_MH_27 0.00988297f
cc_236 N_MM24_g N_MM12_g 0.0171819f
cc_237 N_GCLKN_16 N_MM0_g 0.0253513f
x_PM_ICGx3_ASAP7_75t_R%CLKN VSS N_MM10_g N_MM20_d N_MM21_d N_CLKN_10 N_CLKN_13
+ N_CLKN_18 N_CLKN_3 N_CLKN_15 N_CLKN_12 N_CLKN_1 N_CLKN_11 N_CLKN_17 N_CLKN_14
+ N_CLKN_16 N_CLKN_4 PM_ICGx3_ASAP7_75t_R%CLKN
cc_238 N_CLKN_10 N_CLK_21 0.000185119f
cc_239 N_CLKN_13 N_CLK_21 0.000185189f
cc_240 N_CLKN_18 N_CLK_20 0.000263922f
cc_241 N_CLKN_3 N_CLK_16 0.000285932f
cc_242 N_CLKN_15 N_CLK_15 0.000293691f
cc_243 N_CLKN_12 N_CLK_15 0.00409448f
cc_244 N_CLKN_1 N_CLK_8 0.000315533f
cc_245 N_CLKN_13 N_CLK_16 0.00501337f
cc_246 N_CLKN_1 N_CLK_1 0.0015249f
cc_247 N_CLKN_11 N_MM21_g 0.0157643f
cc_248 N_CLKN_17 N_CLK_17 0.000474087f
cc_249 N_CLKN_15 N_CLK_23 0.000516958f
cc_250 N_CLKN_13 N_CLK_23 0.000698225f
cc_251 N_CLKN_14 N_CLK_15 0.000832624f
cc_252 N_CLKN_16 N_CLK_16 0.00093557f
cc_253 N_CLKN_3 N_MM21_g 0.00094502f
cc_254 N_CLKN_3 N_CLK_3 0.000965282f
cc_255 N_CLKN_4 N_MM21_g 0.00135352f
cc_256 N_CLKN_1 N_CLK_2 0.00147977f
cc_257 N_MM10_g N_MM1_g 0.00161645f
cc_258 N_CLKN_11 N_CLK_3 0.0016435f
cc_259 N_CLKN_17 N_CLK_21 0.00174329f
cc_260 N_MM10_g N_MM9_g 0.00909952f
cc_261 N_CLKN_18 N_CLK_23 0.0263078f
cc_262 N_CLKN_10 N_MM21_g 0.05417f
x_PM_ICGx3_ASAP7_75t_R%CLK VSS CLK N_MM1_g N_MM9_g N_MM21_g N_MM16_g N_MM13_g
+ N_CLK_23 N_CLK_1 N_CLK_15 N_CLK_21 N_CLK_20 N_CLK_16 N_CLK_8 N_CLK_17 N_CLK_3
+ N_CLK_2 N_CLK_19 N_CLK_22 N_CLK_4 N_CLK_18 PM_ICGx3_ASAP7_75t_R%CLK
cc_263 N_CLK_23 N_NET14_14 0.000618672f
cc_264 N_CLK_1 N_NET14_1 0.00159338f
cc_265 N_MM1_g N_MM3_g 0.00327215f
cc_266 N_CLK_15 N_NET14_14 0.0045983f
*END of ICGx3_ASAP7_75t_R.pxi
.ENDS
** Design:	DHLx1_ASAP7_75t_R
* Created:	"Fri Aug 17 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "DHLx1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "DHLx1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_DHLx1_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.0418707f
.ends

.subckt PM_DHLx1_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.0418263f
.ends

.subckt PM_DHLx1_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.00466808f
.ends

.subckt PM_DHLx1_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.00453021f
.ends

.subckt PM_DHLx1_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.00480381f
.ends

.subckt PM_DHLx1_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.0417615f
.ends

.subckt PM_DHLx1_ASAP7_75t_R%Q VSS 17 13 25 7 11 1 2 8 9
c1 1 VSS 0.00872983f
c2 2 VSS 0.00880902f
c3 7 VSS 0.00374654f
c4 8 VSS 0.00374264f
c5 9 VSS 0.0039192f
c6 10 VSS 0.00647246f
c7 11 VSS 0.00582043f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7415 $Y=0.2025 $X2=0.7540 $Y2=0.2025
r2 25 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.2025 $X2=0.7415 $Y2=0.2025
r3 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7560 $Y=0.2025
+ $X2=0.7560 $Y2=0.2340
r4 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.2340 $X2=0.7695 $Y2=0.2340
r5 11 20 7.6809 $w=1.41842e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7830 $Y=0.2340 $X2=0.7830 $Y2=0.1960
r6 11 23 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7830 $Y=0.2340 $X2=0.7695 $Y2=0.2340
r7 19 20 12.0093 $w=1.3e-08 $l=5.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1445 $X2=0.7830 $Y2=0.1960
r8 18 19 9.96886 $w=1.3e-08 $l=4.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1017 $X2=0.7830 $Y2=0.1445
r9 17 18 4.83869 $w=1.3e-08 $l=2.07e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.0810 $X2=0.7830 $Y2=0.1017
r10 17 9 4.25571 $w=1.3e-08 $l=1.83e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.0810 $X2=0.7830 $Y2=0.0627
r11 9 16 5.05752 $w=1.46822e-08 $l=2.67e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7830 $Y=0.0627 $X2=0.7830 $Y2=0.0360
r12 15 16 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7695 $Y=0.0360 $X2=0.7830 $Y2=0.0360
r13 14 15 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.0360 $X2=0.7695 $Y2=0.0360
r14 10 14 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.7445
+ $Y=0.0360 $X2=0.7560 $Y2=0.0360
r15 1 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7560 $Y=0.0675
+ $X2=0.7560 $Y2=0.0360
r16 7 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7415 $Y=0.0675 $X2=0.7540 $Y2=0.0675
r17 13 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.0675 $X2=0.7415 $Y2=0.0675
.ends

.subckt PM_DHLx1_ASAP7_75t_R%PD3 VSS 2 4 1
c1 1 VSS 0.000885753f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0405 $X2=0.4905 $Y2=0.0405
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0405 $X2=0.4735 $Y2=0.0405
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4735 $Y=0.0405 $X2=0.4905 $Y2=0.0405
.ends

.subckt PM_DHLx1_ASAP7_75t_R%PU1 VSS 2 4 1
c1 1 VSS 0.000958663f
r1 4 3 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3365 $Y2=0.2025
r2 2 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3195 $Y2=0.2025
r3 1 3 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3195 $Y=0.2025 $X2=0.3365 $Y2=0.2025
.ends

.subckt PM_DHLx1_ASAP7_75t_R%PD1 VSS 7 10 5 4 1
c1 1 VSS 0.00958371f
c2 4 VSS 0.00317927f
c3 5 VSS 0.0018775f
r1 10 9 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r2 8 9 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r3 5 8 0.123457 $w=8.1e-08 $l=1e-08 $layer=N_src_drn $thickness=1e-09 $X=0.3780
+ $Y=0.0675 $X2=0.3880 $Y2=0.0675
r4 4 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3220 $Y2=0.0675
r5 7 4 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r6 1 5 1e-05
.ends

.subckt PM_DHLx1_ASAP7_75t_R%CLK VSS 11 3 8 6 1 4 7 5
c1 1 VSS 0.00251916f
c2 3 VSS 0.0596925f
c3 4 VSS 0.000775496f
c4 5 VSS 0.00423071f
c5 6 VSS 0.00410402f
c6 7 VSS 0.0019051f
c7 8 VSS 0.00165612f
r1 6 17 1.35805 $w=2.83333e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.1935 $X2=0.1080 $Y2=0.1710
r2 5 15 4.50612 $w=2.06667e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0630 $X2=0.1080 $Y2=0.0990
r3 16 17 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.1710 $X2=0.1080 $Y2=0.1710
r4 8 13 1.35805 $w=2.83333e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1710 $X2=0.0810 $Y2=0.1485
r5 8 16 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1710 $X2=0.0945 $Y2=0.1710
r6 14 15 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.0990 $X2=0.1080 $Y2=0.0990
r7 7 10 0.483592 $w=3.42308e-08 $l=1.87e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0990 $X2=0.0810 $Y2=0.1177
r8 7 14 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0990 $X2=0.0945 $Y2=0.0990
r9 11 12 0.874462 $w=1.3e-08 $l=3.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1227
r10 11 10 0.291487 $w=1.3e-08 $l=1.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1177
r11 4 12 2.85657 $w=1.3e-08 $l=1.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1227
r12 4 13 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1485
r13 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r14 1 4 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_DHLx1_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00424371f
.ends

.subckt PM_DHLx1_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.00466169f
.ends

.subckt PM_DHLx1_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.00366374f
.ends

.subckt PM_DHLx1_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.0419587f
.ends

.subckt PM_DHLx1_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00422441f
.ends

.subckt PM_DHLx1_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.0046885f
.ends

.subckt PM_DHLx1_ASAP7_75t_R%PD2 VSS 7 13 5 1 4
c1 1 VSS 0.00766681f
c2 4 VSS 0.00187326f
c3 5 VSS 0.00233671f
r1 13 12 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r2 5 12 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4880 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r3 10 5 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4725
+ $Y=0.2295 $X2=0.4860 $Y2=0.2295
r4 9 10 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4590
+ $Y=0.2295 $X2=0.4725 $Y2=0.2295
r5 8 9 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4455
+ $Y=0.2295 $X2=0.4590 $Y2=0.2295
r6 1 8 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4320
+ $Y=0.2295 $X2=0.4455 $Y2=0.2295
r7 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2295 $X2=0.4300 $Y2=0.2295
r8 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2295 $X2=0.4175 $Y2=0.2295
.ends

.subckt PM_DHLx1_ASAP7_75t_R%D VSS 9 3 4 1 5
c1 1 VSS 0.00720719f
c2 3 VSS 0.0839248f
c3 4 VSS 0.00888442f
c4 5 VSS 0.0071517f
r1 10 11 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1215 $X2=0.2970 $Y2=0.1350
r2 9 10 1.16595 $w=1.3e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1165 $X2=0.2970 $Y2=0.1215
r3 9 8 1.28254 $w=1.3e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1165 $X2=0.2970 $Y2=0.1110
r4 4 8 8.27824 $w=1.3e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0755 $X2=0.2970 $Y2=0.1110
r5 4 5 8.03069 $w=1.41392e-08 $l=3.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0755 $X2=0.2970 $Y2=0.0360
r6 3 1 6.51726 $w=1.18568e-07 $l=5e-10 $layer=LIG $thickness=5.19024e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2970 $Y2=0.1345
r7 1 11 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1345
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_DHLx1_ASAP7_75t_R%NET088 VSS 9 35 41 11 16 1 4 14 3 13 15 10 12
c1 1 VSS 0.00291481f
c2 3 VSS 0.00605459f
c3 4 VSS 0.00643231f
c4 9 VSS 0.0375418f
c5 10 VSS 0.00345804f
c6 11 VSS 0.00363842f
c7 12 VSS 0.00125523f
c8 13 VSS 0.0085738f
c9 14 VSS 0.00557943f
c10 15 VSS 0.00281862f
c11 16 VSS 0.00597496f
c12 17 VSS 0.00369672f
r1 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2295 $X2=0.5920 $Y2=0.2295
r2 41 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.2295 $X2=0.5795 $Y2=0.2295
r3 4 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2295
+ $X2=0.5940 $Y2=0.2340
r4 37 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.2340 $X2=0.6075 $Y2=0.2340
r5 16 33 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.2340 $X2=0.6210 $Y2=0.2160
r6 16 38 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.2340 $X2=0.6075 $Y2=0.2340
r7 10 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.0405 $X2=0.5920 $Y2=0.0405
r8 35 10 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0405 $X2=0.5795 $Y2=0.0405
r9 32 33 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1870 $X2=0.6210 $Y2=0.2160
r10 31 32 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1655 $X2=0.6210 $Y2=0.1870
r11 30 31 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1515 $X2=0.6210 $Y2=0.1655
r12 29 30 4.89699 $w=1.3e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1305 $X2=0.6210 $Y2=0.1515
r13 28 29 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1215 $X2=0.6210 $Y2=0.1305
r14 27 28 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1085 $X2=0.6210 $Y2=0.1215
r15 14 17 6.39593 $w=1.55565e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.0705 $X2=0.6210 $Y2=0.0360
r16 14 27 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0705 $X2=0.6210 $Y2=0.1085
r17 3 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0405
+ $X2=0.5940 $Y2=0.0360
r18 17 26 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.0360 $X2=0.6075 $Y2=0.0360
r19 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0360 $X2=0.6075 $Y2=0.0360
r20 24 25 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5830
+ $Y=0.0360 $X2=0.5940 $Y2=0.0360
r21 13 15 7.32869 $w=1.41688e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5515 $Y=0.0360 $X2=0.5130 $Y2=0.0360
r22 13 24 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5515
+ $Y=0.0360 $X2=0.5830 $Y2=0.0360
r23 12 22 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0590 $X2=0.5130 $Y2=0.0820
r24 12 15 3.71425 $w=1.68348e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.0590 $X2=0.5130 $Y2=0.0360
r25 1 19 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.5130
+ $Y=0.0820 $X2=0.5130 $Y2=0.0820
r26 1 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.0820
+ $X2=0.5130 $Y2=0.0820
r27 9 19 0.314665 $w=2.27e-07 $l=5.3e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5130 $Y2=0.0820
.ends

.subckt PM_DHLx1_ASAP7_75t_R%CLKN VSS 14 15 16 99 101 31 24 28 30 7 6 17 18 1
+ 22 19 23 33 21 32 2 25 8 3 26 27 29 20
c1 1 VSS 0.0016564f
c2 2 VSS 0.000291703f
c3 3 VSS 8.65215e-20
c4 6 VSS 0.00769981f
c5 7 VSS 0.00753626f
c6 8 VSS 0.00483305f
c7 14 VSS 0.0594349f
c8 15 VSS 0.00569284f
c9 16 VSS 0.00508656f
c10 17 VSS 0.00587503f
c11 18 VSS 0.00588081f
c12 19 VSS 0.00688185f
c13 20 VSS 0.0015615f
c14 21 VSS 0.00478411f
c15 22 VSS 0.00374675f
c16 23 VSS 0.000520311f
c17 24 VSS 0.000258515f
c18 25 VSS 0.00092161f
c19 26 VSS 0.00159419f
c20 27 VSS 0.00359811f
c21 28 VSS 0.00159916f
c22 29 VSS 0.00372944f
c23 30 VSS 0.000798692f
c24 31 VSS 0.000415145f
c25 32 VSS 0.000626818f
c26 33 VSS 0.0198094f
r1 14 93 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1340 $Y2=0.1350
r2 101 100 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r3 18 100 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r4 99 98 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r5 17 98 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r6 93 94 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.1340
+ $Y=0.1350 $X2=0.1440 $Y2=0.1350
r7 1 94 1.73797 $w=1.72143e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1475 $Y=0.1350 $X2=0.1440 $Y2=0.1350
r8 1 96 4.72579 $w=1.53e-08 $l=8e-09 $layer=LIG $thickness=4.8e-08 $X=0.1475
+ $Y=0.1350 $X2=0.1555 $Y2=0.1350
r9 7 87 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0550 $Y2=0.2340
r10 6 84 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0550 $Y2=0.0360
r11 23 89 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.1545
+ $Y=0.1350 $X2=0.1705 $Y2=0.1350
r12 23 96 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1545 $Y=0.1350
+ $X2=0.1555 $Y2=0.1350
r13 86 87 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.2340 $X2=0.0550 $Y2=0.2340
r14 22 86 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0460 $Y2=0.2340
r15 22 29 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0180 $Y2=0.2340
r16 83 84 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.0360 $X2=0.0550 $Y2=0.0360
r17 21 83 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0460 $Y2=0.0360
r18 21 27 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0180 $Y2=0.0360
r19 3 73 5.67512 $w=2.4e-08 $l=5e-09 $layer=LISD $thickness=4.02632e-08
+ $X=0.4590 $Y=0.1790 $X2=0.4640 $Y2=0.1790
r20 16 3 2.88446 $w=1.16273e-07 $l=4.4e-08 $layer=LIG $thickness=5.16364e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4590 $Y2=0.1790
r21 31 67 1.49895 $w=1.95333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1890 $Y2=0.1485
r22 31 89 2.6649 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1705 $Y2=0.1350
r23 27 66 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.0360 $X2=0.0180 $Y2=0.0630
r24 71 73 11.0623 $w=2.14976e-08 $l=2.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4845 $Y=0.1790 $X2=0.4640 $Y2=0.1790
r25 70 71 8.84105 $w=2.02e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4995 $Y=0.1790 $X2=0.4845 $Y2=0.1790
r26 8 68 6.18874 $w=2.02e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5025 $Y=0.1790 $X2=0.5130 $Y2=0.1790
r27 8 70 1.76821 $w=2.02e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.5025
+ $Y=0.1790 $X2=0.4995 $Y2=0.1790
r28 24 61 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1665 $X2=0.1890 $Y2=0.1890
r29 24 67 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1665 $X2=0.1890 $Y2=0.1485
r30 20 28 3.9134 $w=1.47857e-08 $l=2.25499e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.2115 $X2=0.0165 $Y2=0.1890
r31 20 29 3.59766 $w=1.692e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.2115 $X2=0.0180 $Y2=0.2340
r32 65 66 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0990 $X2=0.0180 $Y2=0.0630
r33 64 65 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1350 $X2=0.0180 $Y2=0.0990
r34 19 28 3.9134 $w=1.47857e-08 $l=2.25499e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1665 $X2=0.0165 $Y2=0.1890
r35 19 64 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1665 $X2=0.0180 $Y2=0.1350
r36 62 68 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5130 $Y=0.1845
+ $X2=0.5130 $Y2=0.1790
r37 26 62 3.96423 $w=1.3e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1675 $X2=0.5130 $Y2=0.1845
r38 60 61 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1755 $Y=0.1890 $X2=0.1890 $Y2=0.1890
r39 59 60 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.1890 $X2=0.1755 $Y2=0.1890
r40 30 59 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1505
+ $Y=0.1890 $X2=0.1620 $Y2=0.1890
r41 56 57 1.90199 $w=1.38333e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.0255 $Y=0.1890 $X2=0.0345 $Y2=0.1890
r42 28 56 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0165
+ $Y=0.1890 $X2=0.0255 $Y2=0.1890
r43 54 62 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.5130 $Y=0.1890
+ $X2=0.5130 $Y2=0.1845
r44 53 54 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.4770
+ $Y=0.1890 $X2=0.5130 $Y2=0.1890
r45 52 53 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M2 $thickness=3.6e-08 $X=0.4320
+ $Y=0.1890 $X2=0.4770 $Y2=0.1890
r46 50 51 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.1620
+ $Y=0.1890 $X2=0.2000 $Y2=0.1890
r47 50 59 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1620 $Y=0.1890
+ $X2=0.1620 $Y2=0.1890
r48 49 50 15.0407 $w=1.3e-08 $l=6.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.0975
+ $Y=0.1890 $X2=0.1620 $Y2=0.1890
r49 48 49 15.0407 $w=1.3e-08 $l=6.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.0330
+ $Y=0.1890 $X2=0.0975 $Y2=0.1890
r50 48 57 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.0330 $Y=0.1890
+ $X2=0.0345 $Y2=0.1890
r51 46 52 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M2 $thickness=3.6e-08 $X=0.3870
+ $Y=0.1890 $X2=0.4320 $Y2=0.1890
r52 45 46 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1890 $X2=0.3870 $Y2=0.1890
r53 33 45 15.2739 $w=1.3e-08 $l=6.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.2855
+ $Y=0.1890 $X2=0.3510 $Y2=0.1890
r54 33 51 19.9377 $w=1.3e-08 $l=8.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.2855
+ $Y=0.1890 $X2=0.2000 $Y2=0.1890
r55 32 42 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.1980 $X2=0.3510 $Y2=0.1845
r56 32 45 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.3510 $Y=0.1980 $X2=0.3510
+ $Y2=0.1890
r57 42 45 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.3510 $Y=0.1845 $X2=0.3510
+ $Y2=0.1890
r58 41 42 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1755 $X2=0.3510 $Y2=0.1845
r59 40 41 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1570 $X2=0.3510 $Y2=0.1755
r60 39 40 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1340 $X2=0.3510 $Y2=0.1570
r61 25 39 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1155 $X2=0.3510 $Y2=0.1340
r62 15 2 6.51726 $w=1.18568e-07 $l=5e-10 $layer=LIG $thickness=5.19024e-08
+ $X=0.3510 $Y=0.1350 $X2=0.3510 $Y2=0.1345
r63 2 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1345
+ $X2=0.3510 $Y2=0.1340
r64 7 18 1e-05
r65 6 17 1e-05
.ends

.subckt PM_DHLx1_ASAP7_75t_R%CLKB VSS 9 45 47 3 4 13 12 10 11 18 15 14 1 17 16
c1 1 VSS 9.81183e-20
c2 3 VSS 0.00696746f
c3 4 VSS 0.00720038f
c4 9 VSS 0.00450449f
c5 10 VSS 0.00586114f
c6 11 VSS 0.00581107f
c7 12 VSS 0.00865863f
c8 13 VSS 0.00852857f
c9 14 VSS 0.00617747f
c10 15 VSS 0.00067503f
c11 16 VSS 0.00357053f
c12 17 VSS 0.00295952f
c13 18 VSS 0.00506654f
r1 11 4 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1600 $Y2=0.2160
r2 47 11 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r3 10 3 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1600 $Y2=0.0540
r4 45 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r5 4 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r6 3 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r7 42 43 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1845 $Y2=0.2340
r8 13 17 4.75866 $w=1.41702e-08 $l=2.72259e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.2340 $X2=0.2430 $Y2=0.2305
r9 13 43 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.1845 $Y2=0.2340
r10 39 40 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1845 $Y2=0.0360
r11 12 16 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.0360 $X2=0.2430 $Y2=0.0360
r12 12 40 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.1845 $Y2=0.0360
r13 17 36 3.70931 $w=1.44474e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.2305 $X2=0.2430 $Y2=0.2115
r14 16 34 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0360 $X2=0.2430 $Y2=0.0630
r15 35 36 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1890 $X2=0.2430 $Y2=0.2115
r16 33 34 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0990 $X2=0.2430 $Y2=0.0630
r17 32 33 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1215 $X2=0.2430 $Y2=0.0990
r18 31 35 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1710 $X2=0.2430 $Y2=0.1890
r19 30 31 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1530 $X2=0.2430 $Y2=0.1710
r20 14 30 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1530
r21 14 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1215
r22 28 29 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1530 $X2=0.4050 $Y2=0.1530
r23 27 28 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1530 $X2=0.3240 $Y2=0.1530
r24 27 30 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.2430 $Y=0.1530
+ $X2=0.2430 $Y2=0.1530
r25 18 27 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.2315
+ $Y=0.1530 $X2=0.2430 $Y2=0.1530
r26 25 29 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4050 $Y=0.1530
+ $X2=0.4050 $Y2=0.1530
r27 24 25 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1435 $X2=0.4050 $Y2=0.1530
r28 23 24 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1340 $X2=0.4050 $Y2=0.1435
r29 15 23 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1155 $X2=0.4050 $Y2=0.1340
r30 9 1 5.63117 $w=1.26721e-07 $l=3e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4050 $Y2=0.1320
r31 1 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1320
+ $X2=0.4050 $Y2=0.1340
.ends

.subckt PM_DHLx1_ASAP7_75t_R%MH VSS 11 12 66 70 74 78 13 17 16 14 19 5 15 25 20
+ 1 26 21 6 18 24 22 2 23
c1 1 VSS 0.000401177f
c2 2 VSS 0.00450805f
c3 5 VSS 0.0060327f
c4 6 VSS 0.00502502f
c5 11 VSS 0.0370211f
c6 12 VSS 0.0802285f
c7 13 VSS 0.00300801f
c8 14 VSS 0.000440809f
c9 15 VSS 0.00349942f
c10 16 VSS 0.000426032f
c11 17 VSS 0.00791564f
c12 18 VSS 0.00374978f
c13 19 VSS 0.00108853f
c14 20 VSS 0.000680997f
c15 21 VSS 0.000712266f
c16 22 VSS 0.00225184f
c17 23 VSS 0.00246306f
c18 24 VSS 4.00654e-20
c19 25 VSS 0.00295097f
c20 26 VSS 0.00702828f
r1 78 77 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r2 76 77 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r3 15 76 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3760 $Y=0.2295 $X2=0.3880 $Y2=0.2295
r4 16 15 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2295 $X2=0.3760 $Y2=0.2295
r5 72 73 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r6 74 72 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.1890 $X2=0.3635 $Y2=0.1890
r7 15 73 0.185185 $w=5.4e-08 $l=1e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r8 70 69 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r9 68 69 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4420 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r10 6 68 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4300 $Y=0.0405 $X2=0.4420 $Y2=0.0405
r11 14 6 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0405 $X2=0.4300 $Y2=0.0405
r12 13 6 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0810 $X2=0.4300 $Y2=0.0810
r13 66 13 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0810 $X2=0.4175 $Y2=0.0810
r14 62 15 15.0298 $w=2.02e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.3780 $Y=0.2045 $X2=0.3780 $Y2=0.1790
r15 5 56 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2295
+ $X2=0.3740 $Y2=0.2340
r16 5 62 14.7351 $w=2.02e-08 $l=2.5e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.3780 $Y=0.2295 $X2=0.3780 $Y2=0.2045
r17 2 50 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7290 $Y=0.1360
+ $X2=0.7290 $Y2=0.1445
r18 12 2 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=0.7290
+ $Y=0.1350 $X2=0.7290 $Y2=0.1360
r19 6 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0405
+ $X2=0.4320 $Y2=0.0360
r20 53 54 1.98211 $w=1.3e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3830
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r21 53 56 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3830
+ $Y=0.2340 $X2=0.3740 $Y2=0.2340
r22 52 54 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r23 17 25 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4320 $Y=0.2340 $X2=0.4590 $Y2=0.2340
r24 17 52 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4050 $Y2=0.2340
r25 22 50 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1245 $X2=0.7290 $Y2=0.1445
r26 18 23 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4320 $Y=0.0360 $X2=0.4590 $Y2=0.0360
r27 25 45 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4590 $Y2=0.2160
r28 48 50 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.7290 $Y=0.1530
+ $X2=0.7290 $Y2=0.1445
r29 47 48 24.6015 $w=1.3e-08 $l=1.055e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.6235 $Y=0.1530 $X2=0.7290 $Y2=0.1530
r30 46 47 29.3819 $w=1.3e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.4975
+ $Y=0.1530 $X2=0.6235 $Y2=0.1530
r31 26 46 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M2 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1530 $X2=0.4975 $Y2=0.1530
r32 26 40 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4590 $Y=0.1530
+ $X2=0.4590 $Y2=0.1530
r33 23 39 6.39593 $w=1.55565e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4590 $Y2=0.0705
r34 44 45 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1980 $X2=0.4590 $Y2=0.2160
r35 43 44 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1800 $X2=0.4590 $Y2=0.1980
r36 42 43 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1675 $X2=0.4590 $Y2=0.1800
r37 41 42 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1630 $X2=0.4590 $Y2=0.1675
r38 40 41 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1530 $X2=0.4590 $Y2=0.1630
r39 20 40 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1415 $X2=0.4590 $Y2=0.1530
r40 20 24 1.50137 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1415 $X2=0.4590 $Y2=0.1300
r41 38 39 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1010 $X2=0.4590 $Y2=0.0705
r42 19 24 2.66732 $w=1.57273e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1135 $X2=0.4590 $Y2=0.1300
r43 19 38 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1135 $X2=0.4590 $Y2=0.1010
r44 24 36 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1300 $X2=0.4860 $Y2=0.1300
r45 35 36 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1300 $X2=0.4860 $Y2=0.1300
r46 21 33 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1300 $X2=0.5670 $Y2=0.1300
r47 21 35 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1300 $X2=0.5130 $Y2=0.1300
r48 32 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1330
+ $X2=0.5670 $Y2=0.1300
r49 1 30 0.590723 $w=1.53e-08 $l=6e-09 $layer=LIG $thickness=4.8e-08 $X=0.5670
+ $Y=0.1240 $X2=0.5670 $Y2=0.1300
r50 1 31 1.77217 $w=1.53e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08 $X=0.5670
+ $Y=0.1240 $X2=0.5670 $Y2=0.1210
r51 30 31 1.18145 $w=1.53e-08 $l=9e-09 $layer=LIG $thickness=4.8e-08 $X=0.5670
+ $Y=0.1300 $X2=0.5670 $Y2=0.1210
r52 30 32 4.72579 $w=1.53e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08 $X=0.5670
+ $Y=0.1300 $X2=0.5670 $Y2=0.1330
r53 11 30 0.314665 $w=2.27e-07 $l=5e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5670 $Y=0.1350 $X2=0.5670 $Y2=0.1300
.ends


*
.SUBCKT DHLx1_ASAP7_75t_R VSS VDD CLK D Q
*
* VSS VSS
* VDD VDD
* CLK CLK
* D D
* Q Q
*
*

MM0 N_MM0_d N_MM0_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2 N_MM2_d N_MM2_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM10_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM6 N_MM6_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM24 N_MM24_d N_MM25_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM12 N_MM12_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM13 N_MM13_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM25 N_MM25_d N_MM25_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "DHLx1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "DHLx1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_DHLx1_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_DHLx1_ASAP7_75t_R%noxref_19
cc_1 N_noxref_19_1 N_MM3_g 0.00136823f
cc_2 N_noxref_19_1 N_CLKB_11 0.000754168f
cc_3 N_noxref_19_1 N_noxref_16_1 0.000465318f
cc_4 N_noxref_19_1 N_noxref_17_1 0.0076963f
cc_5 N_noxref_19_1 N_noxref_18_1 0.0012342f
x_PM_DHLx1_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_DHLx1_ASAP7_75t_R%noxref_18
cc_6 N_noxref_18_1 N_MM3_g 0.00136072f
cc_7 N_noxref_18_1 N_CLKB_10 0.000788721f
cc_8 N_noxref_18_1 N_noxref_16_1 0.00769881f
cc_9 N_noxref_18_1 N_noxref_17_1 0.000464979f
x_PM_DHLx1_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_DHLx1_ASAP7_75t_R%noxref_20
cc_10 N_noxref_20_1 N_NET088_10 0.0169636f
cc_11 N_noxref_20_1 N_MM7_g 0.00586117f
x_PM_DHLx1_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_DHLx1_ASAP7_75t_R%noxref_25
cc_12 N_noxref_25_1 N_MM25_g 0.00148587f
cc_13 N_noxref_25_1 N_Q_8 0.038586f
cc_14 N_noxref_25_1 N_noxref_24_1 0.00177936f
x_PM_DHLx1_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_DHLx1_ASAP7_75t_R%noxref_24
cc_15 N_noxref_24_1 N_MM25_g 0.00148555f
cc_16 N_noxref_24_1 N_Q_7 0.0383821f
x_PM_DHLx1_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_DHLx1_ASAP7_75t_R%noxref_22
cc_17 N_noxref_22_1 N_NET088_10 0.000560604f
cc_18 N_noxref_22_1 N_MM25_g 0.0016195f
cc_19 N_noxref_22_1 N_noxref_20_1 0.00775007f
cc_20 N_noxref_22_1 N_noxref_21_1 0.000449852f
x_PM_DHLx1_ASAP7_75t_R%Q VSS Q N_MM24_d N_MM25_d N_Q_7 N_Q_11 N_Q_1 N_Q_2 N_Q_8
+ N_Q_9 PM_DHLx1_ASAP7_75t_R%Q
cc_21 N_Q_7 N_MH_22 0.000768093f
cc_22 N_Q_7 N_MH_2 0.000921277f
cc_23 N_Q_11 N_MH_26 0.000978373f
cc_24 N_Q_1 N_MM25_g 0.00107376f
cc_25 N_Q_2 N_MM25_g 0.00119492f
cc_26 N_Q_8 N_MH_2 0.00170812f
cc_27 N_Q_9 N_MH_22 0.00427544f
cc_28 N_Q_8 N_MM25_g 0.0154728f
cc_29 N_Q_7 N_MM25_g 0.0545414f
x_PM_DHLx1_ASAP7_75t_R%PD3 VSS N_MM9_s N_MM8_d N_PD3_1 PM_DHLx1_ASAP7_75t_R%PD3
cc_30 N_PD3_1 N_MM9_g 0.00773043f
cc_31 N_PD3_1 N_MM11_g 0.00779705f
x_PM_DHLx1_ASAP7_75t_R%PU1 VSS N_MM3_d N_MM1_s N_PU1_1 PM_DHLx1_ASAP7_75t_R%PU1
cc_32 N_PU1_1 N_MM1_g 0.0170767f
cc_33 N_PU1_1 N_MM3_g 0.0170358f
x_PM_DHLx1_ASAP7_75t_R%PD1 VSS N_MM5_d N_MM4_s N_PD1_5 N_PD1_4 N_PD1_1
+ PM_DHLx1_ASAP7_75t_R%PD1
cc_34 N_PD1_5 N_CLKN_25 0.000461481f
cc_35 N_PD1_5 N_CLKN_2 0.0024966f
cc_36 N_PD1_5 N_MM1_g 0.0737354f
cc_37 N_PD1_4 N_D_1 0.000644331f
cc_38 N_PD1_4 N_D_4 0.000738572f
cc_39 N_PD1_4 N_MM3_g 0.036113f
cc_40 N_PD1_5 N_CLKB_1 0.000659826f
cc_41 N_PD1_5 N_MM10_g 0.0347944f
cc_42 N_PD1_1 N_MH_18 0.000163069f
cc_43 N_PD1_1 N_MH_6 0.00139658f
cc_44 N_PD1_1 N_MH_13 0.00319858f
x_PM_DHLx1_ASAP7_75t_R%CLK VSS CLK N_MM0_g N_CLK_8 N_CLK_6 N_CLK_1 N_CLK_4
+ N_CLK_7 N_CLK_5 PM_DHLx1_ASAP7_75t_R%CLK
x_PM_DHLx1_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_DHLx1_ASAP7_75t_R%noxref_15
cc_45 N_noxref_15_1 N_MM0_g 0.00367732f
cc_46 N_noxref_15_1 N_CLKN_29 5.45631e-20
cc_47 N_noxref_15_1 N_CLKN_20 8.02427e-20
cc_48 N_noxref_15_1 N_CLKN_28 8.9607e-20
cc_49 N_noxref_15_1 N_CLKN_19 0.000271578f
cc_50 N_noxref_15_1 N_CLKN_7 0.000435397f
cc_51 N_noxref_15_1 N_CLKN_18 0.0277721f
cc_52 N_noxref_15_1 N_noxref_14_1 0.00204815f
x_PM_DHLx1_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_DHLx1_ASAP7_75t_R%noxref_17
cc_53 N_noxref_17_1 N_CLKN_1 0.000395083f
cc_54 N_noxref_17_1 N_MM2_g 0.00366263f
cc_55 N_noxref_17_1 N_CLKB_11 0.0274329f
cc_56 N_noxref_17_1 N_noxref_16_1 0.00141536f
x_PM_DHLx1_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_DHLx1_ASAP7_75t_R%noxref_21
cc_57 N_noxref_21_1 N_CLKN_8 0.00288986f
cc_58 N_noxref_21_1 N_NET088_11 0.0163772f
cc_59 N_noxref_21_1 N_MM7_g 0.00527943f
cc_60 N_noxref_21_1 N_noxref_20_1 0.00148426f
x_PM_DHLx1_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_DHLx1_ASAP7_75t_R%noxref_23
cc_61 N_noxref_23_1 N_CLKN_8 0.000605158f
cc_62 N_noxref_23_1 N_MM25_g 0.00156599f
cc_63 N_noxref_23_1 N_noxref_20_1 0.000470346f
cc_64 N_noxref_23_1 N_noxref_21_1 0.00760963f
cc_65 N_noxref_23_1 N_noxref_22_1 0.00122905f
x_PM_DHLx1_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_DHLx1_ASAP7_75t_R%noxref_14
cc_66 N_noxref_14_1 N_MM0_g 0.00370893f
cc_67 N_noxref_14_1 N_CLKN_6 0.00048495f
cc_68 N_noxref_14_1 N_CLKN_27 5.92385e-20
cc_69 N_noxref_14_1 N_CLKN_19 0.000382798f
cc_70 N_noxref_14_1 N_CLKN_17 0.0276706f
x_PM_DHLx1_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_DHLx1_ASAP7_75t_R%noxref_16
cc_71 N_noxref_16_1 N_CLKN_1 0.00039096f
cc_72 N_noxref_16_1 N_MM2_g 0.00357605f
cc_73 N_noxref_16_1 N_CLKB_10 0.0274831f
x_PM_DHLx1_ASAP7_75t_R%PD2 VSS N_MM10_s N_MM11_d N_PD2_5 N_PD2_1 N_PD2_4
+ PM_DHLx1_ASAP7_75t_R%PD2
cc_74 N_PD2_5 N_CLKN_8 0.00125881f
cc_75 N_PD2_1 N_CLKN_3 0.000886031f
cc_76 N_PD2_1 N_MM9_g 0.00219475f
cc_77 N_PD2_4 N_MM9_g 0.0071504f
cc_78 N_PD2_5 N_MM9_g 0.0240485f
cc_79 N_PD2_4 N_MM10_g 0.0150536f
cc_80 N_PD2_5 N_MM11_g 0.0146108f
cc_81 N_PD2_1 N_MH_15 0.000618569f
cc_82 N_PD2_1 N_MH_17 0.000420174f
cc_83 N_PD2_1 N_MH_20 0.000432258f
cc_84 N_PD2_4 N_MH_5 0.000615419f
cc_85 N_PD2_1 N_MH_25 0.0021199f
x_PM_DHLx1_ASAP7_75t_R%D VSS D N_MM3_g N_D_4 N_D_1 N_D_5 PM_DHLx1_ASAP7_75t_R%D
cc_86 N_D_4 N_CLKN_32 0.000573213f
cc_87 N_D_4 N_CLKN_33 0.000833394f
cc_88 N_D_1 N_CLKN_2 0.0023237f
cc_89 N_MM3_g N_MM1_g 0.00506514f
cc_90 N_D_4 N_CLKN_25 0.00554127f
x_PM_DHLx1_ASAP7_75t_R%NET088 VSS N_MM11_g N_MM6_d N_MM7_d N_NET088_11
+ N_NET088_16 N_NET088_1 N_NET088_4 N_NET088_14 N_NET088_3 N_NET088_13
+ N_NET088_15 N_NET088_10 N_NET088_12 PM_DHLx1_ASAP7_75t_R%NET088
cc_91 N_MM11_g N_CLKN_26 0.000371837f
cc_92 N_MM11_g N_CLKN_8 0.00513228f
cc_93 N_MM11_g N_CLKN_3 0.000148702f
cc_94 N_MM11_g N_CLKN_33 0.000192524f
cc_95 N_NET088_11 N_CLKN_8 0.00038882f
cc_96 N_NET088_16 N_CLKN_8 0.000414286f
cc_97 N_NET088_1 N_MM9_g 0.00042377f
cc_98 N_NET088_4 N_CLKN_8 0.000892611f
cc_99 N_NET088_14 N_CLKN_8 0.00135816f
cc_100 N_MM11_g N_MM9_g 0.0143353f
x_PM_DHLx1_ASAP7_75t_R%CLKN VSS N_MM2_g N_MM1_g N_MM9_g N_MM0_d N_MM12_d
+ N_CLKN_31 N_CLKN_24 N_CLKN_28 N_CLKN_30 N_CLKN_7 N_CLKN_6 N_CLKN_17 N_CLKN_18
+ N_CLKN_1 N_CLKN_22 N_CLKN_19 N_CLKN_23 N_CLKN_33 N_CLKN_21 N_CLKN_32 N_CLKN_2
+ N_CLKN_25 N_CLKN_8 N_CLKN_3 N_CLKN_26 N_CLKN_27 N_CLKN_29 N_CLKN_20
+ PM_DHLx1_ASAP7_75t_R%CLKN
cc_101 N_CLKN_31 N_MM0_g 7.58761e-20
cc_102 N_CLKN_24 N_MM0_g 0.000107013f
cc_103 N_CLKN_28 N_MM0_g 0.000184101f
cc_104 N_CLKN_30 N_MM0_g 0.000187475f
cc_105 N_CLKN_7 N_MM0_g 0.00107419f
cc_106 N_CLKN_6 N_MM0_g 0.00115113f
cc_107 N_CLKN_17 N_MM0_g 0.0112216f
cc_108 N_CLKN_18 N_MM0_g 0.0113259f
cc_109 N_CLKN_1 N_CLK_8 0.000441107f
cc_110 N_CLKN_22 N_CLK_6 0.000655904f
cc_111 N_CLKN_1 N_CLK_1 0.00331106f
cc_112 N_CLKN_19 N_CLK_4 0.00106325f
cc_113 N_CLKN_23 N_CLK_8 0.00120365f
cc_114 N_CLKN_23 N_CLK_7 0.00139667f
cc_115 N_CLKN_33 N_CLK_8 0.00164872f
cc_116 N_CLKN_30 N_CLK_6 0.00168087f
cc_117 N_CLKN_21 N_CLK_5 0.001733f
cc_118 N_CLKN_30 N_CLK_8 0.00219674f
cc_119 N_CLKN_28 N_CLK_8 0.0029115f
cc_120 N_CLKN_19 N_CLK_7 0.0029493f
cc_121 N_MM2_g N_MM0_g 0.0351454f
x_PM_DHLx1_ASAP7_75t_R%CLKB VSS N_MM10_g N_MM2_d N_MM13_d N_CLKB_3 N_CLKB_4
+ N_CLKB_13 N_CLKB_12 N_CLKB_10 N_CLKB_11 N_CLKB_18 N_CLKB_15 N_CLKB_14
+ N_CLKB_1 N_CLKB_17 N_CLKB_16 PM_DHLx1_ASAP7_75t_R%CLKB
cc_122 N_CLKB_3 N_CLK_5 0.000437879f
cc_123 N_CLKB_4 N_CLK_5 0.00019816f
cc_124 N_CLKB_13 N_CLK_6 0.00106614f
cc_125 N_CLKB_12 N_CLK_5 0.00274652f
cc_126 N_CLKB_10 N_CLKN_19 5.8821e-20
cc_127 N_CLKB_10 N_CLKN_8 0.000115256f
cc_128 N_CLKB_10 N_CLKN_30 0.000221545f
cc_129 N_CLKB_4 N_CLKN_30 0.000283373f
cc_130 N_CLKB_13 N_CLKN_30 0.00474673f
cc_131 N_CLKB_11 N_MM2_g 0.0111457f
cc_132 N_CLKB_18 N_CLKN_25 0.000395204f
cc_133 N_CLKB_4 N_CLKN_1 0.000415101f
cc_134 N_CLKB_12 N_CLKN_31 0.0004488f
cc_135 N_CLKB_15 N_CLKN_32 0.000492957f
cc_136 N_CLKB_14 N_CLKN_23 0.000601159f
cc_137 N_CLKB_15 N_CLKN_33 0.000665257f
cc_138 N_MM10_g N_CLKN_3 0.000675128f
cc_139 N_CLKB_3 N_MM2_g 0.00074301f
cc_140 N_CLKB_11 N_CLKN_1 0.000901256f
cc_141 N_CLKB_1 N_CLKN_2 0.00226448f
cc_142 N_CLKB_14 N_CLKN_33 0.000938226f
cc_143 N_CLKB_4 N_MM2_g 0.00111127f
cc_144 N_CLKB_14 N_CLKN_24 0.0011563f
cc_145 N_MM10_g N_MM1_g 0.00162868f
cc_146 N_CLKB_14 N_CLKN_31 0.00377864f
cc_147 N_CLKB_15 N_CLKN_25 0.00386238f
cc_148 N_MM10_g N_MM9_g 0.00909008f
cc_149 N_CLKB_18 N_CLKN_33 0.0186216f
cc_150 N_CLKB_10 N_MM2_g 0.038936f
cc_151 N_CLKB_17 N_D_4 0.000307404f
cc_152 N_CLKB_16 N_D_5 0.000948602f
cc_153 N_CLKB_18 N_D_4 0.00103782f
cc_154 N_CLKB_14 N_D_4 0.00850275f
x_PM_DHLx1_ASAP7_75t_R%MH VSS N_MM7_g N_MM25_g N_MM4_d N_MM9_d N_MM1_d N_MM10_d
+ N_MH_13 N_MH_17 N_MH_16 N_MH_14 N_MH_19 N_MH_5 N_MH_15 N_MH_25 N_MH_20 N_MH_1
+ N_MH_26 N_MH_21 N_MH_6 N_MH_18 N_MH_24 N_MH_22 N_MH_2 N_MH_23
+ PM_DHLx1_ASAP7_75t_R%MH
cc_155 N_MH_13 N_CLKN_26 0.000124991f
cc_156 N_MH_17 N_CLKN_25 0.000132722f
cc_157 N_MH_16 N_MM1_g 0.000151732f
cc_158 N_MH_14 N_MM9_g 0.000170254f
cc_159 N_MH_19 N_CLKN_26 0.000243187f
cc_160 N_MH_5 N_CLKN_2 0.000250516f
cc_161 N_MH_15 N_MM1_g 0.0346148f
cc_162 N_MH_5 N_CLKN_32 0.000312376f
cc_163 N_MH_25 N_CLKN_26 0.000411728f
cc_164 N_MH_20 N_CLKN_33 0.000468675f
cc_165 N_MH_5 N_CLKN_25 0.000525484f
cc_166 N_MH_1 N_CLKN_8 0.00175357f
cc_167 N_MH_26 N_CLKN_26 0.000650185f
cc_168 N_MH_21 N_CLKN_8 0.000651709f
cc_169 N_MH_6 N_MM9_g 0.000660894f
cc_170 N_MH_15 N_CLKN_2 0.000774744f
cc_171 N_MH_20 N_CLKN_3 0.000929711f
cc_172 N_MH_5 N_MM1_g 0.00194946f
cc_173 N_MH_21 N_CLKN_26 0.00199274f
cc_174 N_MH_17 N_CLKN_32 0.00364442f
cc_175 N_MH_26 N_CLKN_33 0.00441619f
cc_176 N_MH_20 N_CLKN_26 0.00460911f
cc_177 N_MH_17 N_CLKN_33 0.00556074f
cc_178 N_MM7_g N_CLKN_8 0.00630582f
cc_179 N_MH_13 N_MM9_g 0.0370284f
cc_180 N_MH_14 N_MM10_g 0.000138687f
cc_181 N_MH_16 N_MM10_g 0.000177764f
cc_182 N_MH_18 N_CLKB_15 0.000245663f
cc_183 N_MH_17 N_CLKB_15 0.000297518f
cc_184 N_MH_15 N_MM10_g 0.0167631f
cc_185 N_MH_26 N_CLKB_18 0.00063966f
cc_186 N_MH_20 N_CLKB_15 0.00176797f
cc_187 N_MH_19 N_CLKB_15 0.000852771f
cc_188 N_MH_6 N_CLKB_1 0.000896545f
cc_189 N_MH_17 N_CLKB_18 0.000902973f
cc_190 N_MH_6 N_MM10_g 0.0011185f
cc_191 N_MH_5 N_MM10_g 0.00118512f
cc_192 N_MH_13 N_CLKB_1 0.00170397f
cc_193 N_MH_24 N_CLKB_15 0.00297933f
cc_194 N_MH_13 N_MM10_g 0.0537765f
cc_195 N_MH_22 N_MM11_g 8.99381e-20
cc_196 N_MH_2 N_MM11_g 9.94854e-20
cc_197 N_MH_13 N_MM11_g 0.000168632f
cc_198 N_MH_21 N_MM11_g 0.000170859f
cc_199 N_MH_22 N_NET088_14 0.000305825f
cc_200 N_MM7_g N_NET088_3 0.000363693f
cc_201 N_MH_26 N_NET088_16 0.000416967f
cc_202 N_MH_6 N_NET088_1 0.000438812f
cc_203 N_MH_21 N_NET088_13 0.000634958f
cc_204 N_MH_1 N_NET088_14 0.000798657f
cc_205 N_MH_23 N_NET088_15 0.000912245f
cc_206 N_MH_21 N_NET088_1 0.000923139f
cc_207 N_MH_1 N_MM11_g 0.000927389f
cc_208 N_MM7_g N_NET088_1 0.00108474f
cc_209 N_MM7_g N_NET088_10 0.00660729f
cc_210 N_MM7_g N_NET088_11 0.00653611f
cc_211 N_MH_26 N_NET088_14 0.00264593f
cc_212 N_MH_21 N_NET088_12 0.00288653f
cc_213 N_MH_19 N_NET088_12 0.00355166f
cc_214 N_MH_21 N_NET088_14 0.00410472f
cc_215 N_MM7_g N_MM11_g 0.02941f
*END of DHLx1_ASAP7_75t_R.pxi
.ENDS
** Design:	DHLx2_ASAP7_75t_R
* Created:	"Fri Aug 17 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "DHLx2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "DHLx2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_DHLx2_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.0418707f
.ends

.subckt PM_DHLx2_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.0418263f
.ends

.subckt PM_DHLx2_ASAP7_75t_R%PU1 VSS 2 4 1
c1 1 VSS 0.000958613f
r1 4 3 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3365 $Y2=0.2025
r2 2 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3195 $Y2=0.2025
r3 1 3 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3195 $Y=0.2025 $X2=0.3365 $Y2=0.2025
.ends

.subckt PM_DHLx2_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00424697f
.ends

.subckt PM_DHLx2_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.00466718f
.ends

.subckt PM_DHLx2_ASAP7_75t_R%CLK VSS 11 3 8 6 1 4 7 5
c1 1 VSS 0.00250819f
c2 3 VSS 0.059687f
c3 4 VSS 0.00077001f
c4 5 VSS 0.00422522f
c5 6 VSS 0.00409854f
c6 7 VSS 0.00188318f
c7 8 VSS 0.00165073f
r1 6 17 1.35805 $w=2.83333e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.1935 $X2=0.1080 $Y2=0.1710
r2 5 15 4.50612 $w=2.06667e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0630 $X2=0.1080 $Y2=0.0990
r3 16 17 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.1710 $X2=0.1080 $Y2=0.1710
r4 8 13 1.35805 $w=2.83333e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1710 $X2=0.0810 $Y2=0.1485
r5 8 16 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1710 $X2=0.0945 $Y2=0.1710
r6 14 15 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.0990 $X2=0.1080 $Y2=0.0990
r7 7 10 0.483592 $w=3.42308e-08 $l=1.87e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0990 $X2=0.0810 $Y2=0.1177
r8 7 14 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0990 $X2=0.0945 $Y2=0.0990
r9 11 12 0.874462 $w=1.3e-08 $l=3.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1227
r10 11 10 0.291487 $w=1.3e-08 $l=1.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1177
r11 4 12 2.85657 $w=1.3e-08 $l=1.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1227
r12 4 13 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1485
r13 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r14 1 4 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_DHLx2_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.00468443f
.ends

.subckt PM_DHLx2_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00422572f
.ends

.subckt PM_DHLx2_ASAP7_75t_R%D VSS 9 3 4 1 5
c1 1 VSS 0.00724064f
c2 3 VSS 0.0839415f
c3 4 VSS 0.00890492f
c4 5 VSS 0.00715074f
r1 10 11 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1215 $X2=0.2970 $Y2=0.1350
r2 9 10 1.16595 $w=1.3e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1165 $X2=0.2970 $Y2=0.1215
r3 9 8 1.28254 $w=1.3e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1165 $X2=0.2970 $Y2=0.1110
r4 4 8 8.27824 $w=1.3e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0755 $X2=0.2970 $Y2=0.1110
r5 4 5 8.03069 $w=1.41392e-08 $l=3.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0755 $X2=0.2970 $Y2=0.0360
r6 3 1 6.51726 $w=1.18568e-07 $l=5e-10 $layer=LIG $thickness=5.19024e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2970 $Y2=0.1345
r7 1 11 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1345
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_DHLx2_ASAP7_75t_R%PD3 VSS 2 4 1
c1 1 VSS 0.000878959f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0405 $X2=0.4905 $Y2=0.0405
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0405 $X2=0.4735 $Y2=0.0405
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4735 $Y=0.0405 $X2=0.4905 $Y2=0.0405
.ends

.subckt PM_DHLx2_ASAP7_75t_R%Q VSS 23 16 17 33 34 7 9 1 10 8 2 11
c1 1 VSS 0.00945763f
c2 2 VSS 0.0100144f
c3 7 VSS 0.00461103f
c4 8 VSS 0.00454253f
c5 9 VSS 0.00808066f
c6 10 VSS 0.00798313f
c7 11 VSS 0.00535015f
c8 12 VSS 0.00202562f
c9 13 VSS 0.002154f
r1 34 32 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.2025 $X2=0.7705 $Y2=0.2025
r2 2 32 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7560 $Y=0.2025 $X2=0.7705 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7415 $Y=0.2025 $X2=0.7560 $Y2=0.2025
r4 33 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.2025 $X2=0.7415 $Y2=0.2025
r5 2 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7560 $Y=0.2025
+ $X2=0.7560 $Y2=0.2250
r6 28 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.2250 $X2=0.7695 $Y2=0.2250
r7 26 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.2250 $X2=0.7695 $Y2=0.2250
r8 9 13 5.11339 $w=1.45517e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8120 $Y=0.2250 $X2=0.8410 $Y2=0.2250
r9 9 26 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.8120
+ $Y=0.2250 $X2=0.7830 $Y2=0.2250
r10 13 25 6.16274 $w=1.56328e-08 $l=3.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8410 $Y=0.2250 $X2=0.8410 $Y2=0.1915
r11 24 25 11.6012 $w=1.3e-08 $l=4.98e-08 $layer=M1 $thickness=3.6e-08 $X=0.8410
+ $Y=0.1417 $X2=0.8410 $Y2=0.1915
r12 23 24 6.00464 $w=1.3e-08 $l=2.57e-08 $layer=M1 $thickness=3.6e-08 $X=0.8410
+ $Y=0.1160 $X2=0.8410 $Y2=0.1417
r13 23 22 3.08976 $w=1.3e-08 $l=1.33e-08 $layer=M1 $thickness=3.6e-08 $X=0.8410
+ $Y=0.1160 $X2=0.8410 $Y2=0.1027
r14 11 12 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8410 $Y=0.0720 $X2=0.8410 $Y2=0.0450
r15 11 22 7.17059 $w=1.3e-08 $l=3.07e-08 $layer=M1 $thickness=3.6e-08 $X=0.8410
+ $Y=0.0720 $X2=0.8410 $Y2=0.1027
r16 12 21 5.11339 $w=1.45517e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8410 $Y=0.0450 $X2=0.8120 $Y2=0.0450
r17 20 21 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.0450 $X2=0.8120 $Y2=0.0450
r18 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7695
+ $Y=0.0450 $X2=0.7830 $Y2=0.0450
r19 18 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.0450 $X2=0.7695 $Y2=0.0450
r20 10 18 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.7445
+ $Y=0.0450 $X2=0.7560 $Y2=0.0450
r21 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7560 $Y=0.0675
+ $X2=0.7560 $Y2=0.0450
r22 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.0675 $X2=0.7705 $Y2=0.0675
r23 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7560 $Y=0.0675 $X2=0.7705 $Y2=0.0675
r24 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7415 $Y=0.0675 $X2=0.7560 $Y2=0.0675
r25 16 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.0675 $X2=0.7415 $Y2=0.0675
.ends

.subckt PM_DHLx2_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.00464179f
.ends

.subckt PM_DHLx2_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.00366287f
.ends

.subckt PM_DHLx2_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.041729f
.ends

.subckt PM_DHLx2_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.0422939f
.ends

.subckt PM_DHLx2_ASAP7_75t_R%PD2 VSS 7 13 5 1 4
c1 1 VSS 0.00766612f
c2 4 VSS 0.00187309f
c3 5 VSS 0.0023365f
r1 13 12 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r2 5 12 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4880 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r3 10 5 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4725
+ $Y=0.2295 $X2=0.4860 $Y2=0.2295
r4 9 10 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4590
+ $Y=0.2295 $X2=0.4725 $Y2=0.2295
r5 8 9 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4455
+ $Y=0.2295 $X2=0.4590 $Y2=0.2295
r6 1 8 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4320
+ $Y=0.2295 $X2=0.4455 $Y2=0.2295
r7 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2295 $X2=0.4300 $Y2=0.2295
r8 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2295 $X2=0.4175 $Y2=0.2295
.ends

.subckt PM_DHLx2_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.041941f
.ends

.subckt PM_DHLx2_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.0423773f
.ends

.subckt PM_DHLx2_ASAP7_75t_R%PD1 VSS 7 10 5 4 1
c1 1 VSS 0.00958289f
c2 4 VSS 0.00317903f
c3 5 VSS 0.00187734f
r1 10 9 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r2 8 9 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r3 5 8 0.123457 $w=8.1e-08 $l=1e-08 $layer=N_src_drn $thickness=1e-09 $X=0.3780
+ $Y=0.0675 $X2=0.3880 $Y2=0.0675
r4 4 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3220 $Y2=0.0675
r5 7 4 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r6 1 5 1e-05
.ends

.subckt PM_DHLx2_ASAP7_75t_R%CLKN VSS 14 15 16 99 101 31 24 28 30 7 6 17 18 1
+ 22 19 23 33 21 25 32 2 8 3 26 27 29 20
c1 1 VSS 0.00165572f
c2 2 VSS 0.000290928f
c3 3 VSS 8.61695e-20
c4 6 VSS 0.00768942f
c5 7 VSS 0.0075261f
c6 8 VSS 0.00482577f
c7 14 VSS 0.0594348f
c8 15 VSS 0.00569921f
c9 16 VSS 0.00507917f
c10 17 VSS 0.00582109f
c11 18 VSS 0.00582752f
c12 19 VSS 0.00677478f
c13 20 VSS 0.00154202f
c14 21 VSS 0.00477106f
c15 22 VSS 0.00374509f
c16 23 VSS 0.000518664f
c17 24 VSS 0.000258413f
c18 25 VSS 0.00084809f
c19 26 VSS 0.00159227f
c20 27 VSS 0.00379201f
c21 28 VSS 0.00157744f
c22 29 VSS 0.00371161f
c23 30 VSS 0.000797045f
c24 31 VSS 0.000411925f
c25 32 VSS 0.000626318f
c26 33 VSS 0.0203495f
r1 101 100 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r2 18 100 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r3 99 98 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r4 17 98 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r5 7 96 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0550 $Y2=0.2340
r6 6 93 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0550 $Y2=0.0360
r7 95 96 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.2340 $X2=0.0550 $Y2=0.2340
r8 22 95 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0460 $Y2=0.2340
r9 22 29 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0180 $Y2=0.2340
r10 92 93 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.0360 $X2=0.0550 $Y2=0.0360
r11 21 92 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0460 $Y2=0.0360
r12 21 27 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0180 $Y2=0.0360
r13 3 82 5.67512 $w=2.4e-08 $l=5e-09 $layer=LISD $thickness=4.02632e-08
+ $X=0.4590 $Y=0.1790 $X2=0.4640 $Y2=0.1790
r14 16 3 2.88446 $w=1.16273e-07 $l=4.4e-08 $layer=LIG $thickness=5.16364e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4590 $Y2=0.1790
r15 15 76 6.51726 $w=1.18568e-07 $l=5e-10 $layer=LIG $thickness=5.19024e-08
+ $X=0.3510 $Y=0.1350 $X2=0.3510 $Y2=0.1345
r16 27 75 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.0360 $X2=0.0180 $Y2=0.0630
r17 80 82 11.0623 $w=2.14976e-08 $l=2.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4845 $Y=0.1790 $X2=0.4640 $Y2=0.1790
r18 79 80 8.84105 $w=2.02e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4995 $Y=0.1790 $X2=0.4845 $Y2=0.1790
r19 8 77 6.18874 $w=2.02e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5025 $Y=0.1790 $X2=0.5130 $Y2=0.1790
r20 8 79 1.76821 $w=2.02e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.5025
+ $Y=0.1790 $X2=0.4995 $Y2=0.1790
r21 2 76 6.49795 $w=1.53e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08 $X=0.3510
+ $Y=0.1235 $X2=0.3510 $Y2=0.1345
r22 20 28 3.9134 $w=1.47857e-08 $l=2.25499e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.2115 $X2=0.0165 $Y2=0.1890
r23 20 29 3.59766 $w=1.692e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.2115 $X2=0.0180 $Y2=0.2340
r24 74 75 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0990 $X2=0.0180 $Y2=0.0630
r25 73 74 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1350 $X2=0.0180 $Y2=0.0990
r26 19 28 3.9134 $w=1.47857e-08 $l=2.25499e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1665 $X2=0.0165 $Y2=0.1890
r27 19 73 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1665 $X2=0.0180 $Y2=0.1350
r28 71 77 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5130 $Y=0.1845
+ $X2=0.5130 $Y2=0.1790
r29 26 71 3.96423 $w=1.3e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1675 $X2=0.5130 $Y2=0.1845
r30 32 65 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.1980 $X2=0.3510 $Y2=0.1845
r31 32 56 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.3510 $Y=0.1980 $X2=0.3510
+ $Y2=0.1890
r32 67 68 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1340 $X2=0.3510 $Y2=0.1570
r33 67 76 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1340
+ $X2=0.3510 $Y2=0.1345
r34 25 65 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1755 $X2=0.3510 $Y2=0.1845
r35 25 68 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1755 $X2=0.3510 $Y2=0.1570
r36 62 63 1.90199 $w=1.38333e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.0255 $Y=0.1890 $X2=0.0345 $Y2=0.1890
r37 28 62 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0165
+ $Y=0.1890 $X2=0.0255 $Y2=0.1890
r38 60 71 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.5130 $Y=0.1890
+ $X2=0.5130 $Y2=0.1845
r39 59 60 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.4770
+ $Y=0.1890 $X2=0.5130 $Y2=0.1890
r40 58 59 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M2 $thickness=3.6e-08 $X=0.4320
+ $Y=0.1890 $X2=0.4770 $Y2=0.1890
r41 57 58 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M2 $thickness=3.6e-08 $X=0.3870
+ $Y=0.1890 $X2=0.4320 $Y2=0.1890
r42 56 57 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1890 $X2=0.3870 $Y2=0.1890
r43 56 65 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.3510 $Y=0.1890 $X2=0.3510
+ $Y2=0.1845
r44 55 56 15.2739 $w=1.3e-08 $l=6.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.2855
+ $Y=0.1890 $X2=0.3510 $Y2=0.1890
r45 54 55 19.9377 $w=1.3e-08 $l=8.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.2000
+ $Y=0.1890 $X2=0.2855 $Y2=0.1890
r46 53 54 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.1620
+ $Y=0.1890 $X2=0.2000 $Y2=0.1890
r47 52 53 15.0407 $w=1.3e-08 $l=6.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.0975
+ $Y=0.1890 $X2=0.1620 $Y2=0.1890
r48 51 52 15.0407 $w=1.3e-08 $l=6.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.0330
+ $Y=0.1890 $X2=0.0975 $Y2=0.1890
r49 51 63 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.0330 $Y=0.1890
+ $X2=0.0345 $Y2=0.1890
r50 33 51 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.0215
+ $Y=0.1890 $X2=0.0330 $Y2=0.1890
r51 49 50 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.1890 $X2=0.1755 $Y2=0.1890
r52 49 53 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1620 $Y=0.1890
+ $X2=0.1620 $Y2=0.1890
r53 30 47 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1890 $X2=0.1890 $Y2=0.1665
r54 30 50 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1890 $X2=0.1755 $Y2=0.1890
r55 24 31 1.49895 $w=1.95333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1485 $X2=0.1890 $Y2=0.1350
r56 24 47 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1485 $X2=0.1890 $Y2=0.1665
r57 31 46 2.6649 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1705 $Y2=0.1350
r58 45 46 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.1545
+ $Y=0.1350 $X2=0.1705 $Y2=0.1350
r59 44 45 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1455
+ $Y=0.1350 $X2=0.1545 $Y2=0.1350
r60 23 44 1.16595 $w=1.3e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1405
+ $Y=0.1350 $X2=0.1455 $Y2=0.1350
r61 42 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1555 $Y=0.1350
+ $X2=0.1545 $Y2=0.1350
r62 41 42 4.72579 $w=1.53e-08 $l=8e-09 $layer=LIG $thickness=4.8e-08 $X=0.1475
+ $Y=0.1350 $X2=0.1555 $Y2=0.1350
r63 39 41 1.73797 $w=1.72143e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1440 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r64 1 39 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.1340
+ $Y=0.1350 $X2=0.1440 $Y2=0.1350
r65 14 1 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1340 $Y2=0.1350
r66 14 41 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r67 7 18 1e-05
r68 6 17 1e-05
.ends

.subckt PM_DHLx2_ASAP7_75t_R%NET088 VSS 9 38 44 11 16 1 4 14 3 13 15 10 12
c1 1 VSS 0.00291257f
c2 3 VSS 0.00605266f
c3 4 VSS 0.0064304f
c4 9 VSS 0.0375414f
c5 10 VSS 0.00336995f
c6 11 VSS 0.00355015f
c7 12 VSS 0.00130024f
c8 13 VSS 0.00866507f
c9 14 VSS 0.00507401f
c10 15 VSS 0.00281537f
c11 16 VSS 0.00676256f
c12 17 VSS 0.00309428f
r1 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2295 $X2=0.5920 $Y2=0.2295
r2 44 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.2295 $X2=0.5795 $Y2=0.2295
r3 4 40 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2295
+ $X2=0.5940 $Y2=0.2340
r4 40 41 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.2340 $X2=0.6075 $Y2=0.2340
r5 16 36 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.2340 $X2=0.6210 $Y2=0.2205
r6 16 41 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.2340 $X2=0.6075 $Y2=0.2340
r7 10 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.0405 $X2=0.5920 $Y2=0.0405
r8 38 10 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0405 $X2=0.5795 $Y2=0.0405
r9 35 36 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.2115 $X2=0.6210 $Y2=0.2205
r10 34 35 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1870 $X2=0.6210 $Y2=0.2115
r11 33 34 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1655 $X2=0.6210 $Y2=0.1870
r12 32 33 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1515 $X2=0.6210 $Y2=0.1655
r13 31 32 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1300 $X2=0.6210 $Y2=0.1515
r14 30 31 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1085 $X2=0.6210 $Y2=0.1300
r15 29 30 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0930 $X2=0.6210 $Y2=0.1085
r16 28 29 4.89699 $w=1.3e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0720 $X2=0.6210 $Y2=0.0930
r17 14 27 1.50855 $w=1.55e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0495 $X2=0.6210 $Y2=0.0405
r18 14 28 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0495 $X2=0.6210 $Y2=0.0720
r19 3 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0405
+ $X2=0.5940 $Y2=0.0360
r20 17 26 1.50855 $w=1.55e-08 $l=1.42302e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.0315 $X2=0.6075 $Y2=0.0360
r21 17 27 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0315 $X2=0.6210 $Y2=0.0405
r22 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0360 $X2=0.6075 $Y2=0.0360
r23 24 25 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5830
+ $Y=0.0360 $X2=0.5940 $Y2=0.0360
r24 13 15 7.32869 $w=1.41688e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5515 $Y=0.0360 $X2=0.5130 $Y2=0.0360
r25 13 24 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5515
+ $Y=0.0360 $X2=0.5830 $Y2=0.0360
r26 12 22 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0590 $X2=0.5130 $Y2=0.0820
r27 12 15 3.71425 $w=1.68348e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.0590 $X2=0.5130 $Y2=0.0360
r28 1 19 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.5130
+ $Y=0.0820 $X2=0.5130 $Y2=0.0820
r29 1 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.0820
+ $X2=0.5130 $Y2=0.0820
r30 9 19 0.314665 $w=2.27e-07 $l=5.3e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5130 $Y2=0.0820
.ends

.subckt PM_DHLx2_ASAP7_75t_R%CLKB VSS 9 45 47 3 4 13 12 10 11 18 15 14 1 17 16
c1 1 VSS 9.82572e-20
c2 3 VSS 0.00696762f
c3 4 VSS 0.00720048f
c4 9 VSS 0.00450448f
c5 10 VSS 0.00587727f
c6 11 VSS 0.00582666f
c7 12 VSS 0.0101145f
c8 13 VSS 0.0085304f
c9 14 VSS 0.00617434f
c10 15 VSS 0.000634104f
c11 16 VSS 0.00357102f
c12 17 VSS 0.00295992f
c13 18 VSS 0.00520475f
r1 11 4 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1600 $Y2=0.2160
r2 47 11 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r3 10 3 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1600 $Y2=0.0540
r4 45 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r5 4 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r6 3 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r7 42 43 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1845 $Y2=0.2340
r8 13 17 4.75866 $w=1.41702e-08 $l=2.72259e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.2340 $X2=0.2430 $Y2=0.2305
r9 13 43 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.1845 $Y2=0.2340
r10 39 40 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1845 $Y2=0.0360
r11 12 16 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.0360 $X2=0.2430 $Y2=0.0360
r12 12 40 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.1845 $Y2=0.0360
r13 17 36 3.70931 $w=1.44474e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.2305 $X2=0.2430 $Y2=0.2115
r14 16 34 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0360 $X2=0.2430 $Y2=0.0630
r15 35 36 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1890 $X2=0.2430 $Y2=0.2115
r16 33 34 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0990 $X2=0.2430 $Y2=0.0630
r17 32 33 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1215 $X2=0.2430 $Y2=0.0990
r18 31 35 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1710 $X2=0.2430 $Y2=0.1890
r19 30 31 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1530 $X2=0.2430 $Y2=0.1710
r20 14 30 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1530
r21 14 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1215
r22 28 29 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1530 $X2=0.4050 $Y2=0.1530
r23 27 28 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1530 $X2=0.3240 $Y2=0.1530
r24 27 30 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.2430 $Y=0.1530
+ $X2=0.2430 $Y2=0.1530
r25 18 27 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.2315
+ $Y=0.1530 $X2=0.2430 $Y2=0.1530
r26 25 29 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4050 $Y=0.1530
+ $X2=0.4050 $Y2=0.1530
r27 24 25 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1435 $X2=0.4050 $Y2=0.1530
r28 23 24 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1340 $X2=0.4050 $Y2=0.1435
r29 15 23 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1155 $X2=0.4050 $Y2=0.1340
r30 9 1 5.63117 $w=1.26721e-07 $l=3e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4050 $Y2=0.1320
r31 1 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1320
+ $X2=0.4050 $Y2=0.1340
.ends

.subckt PM_DHLx2_ASAP7_75t_R%MH VSS 13 14 15 77 81 86 90 16 20 19 17 22 7 18 29
+ 23 1 30 24 8 21 28 2 25 27 26 3
c1 1 VSS 0.000424745f
c2 2 VSS 0.00474989f
c3 3 VSS 0.00422542f
c4 7 VSS 0.00605193f
c5 8 VSS 0.00503613f
c6 13 VSS 0.0370215f
c7 14 VSS 0.0803154f
c8 15 VSS 0.0804328f
c9 16 VSS 0.00442649f
c10 17 VSS 0.00110394f
c11 18 VSS 0.00486559f
c12 19 VSS 0.00110222f
c13 20 VSS 0.00818304f
c14 21 VSS 0.0039905f
c15 22 VSS 0.00140084f
c16 23 VSS 0.000694628f
c17 24 VSS 0.000558852f
c18 25 VSS 0.00346713f
c19 26 VSS 0.0028103f
c20 27 VSS 0.00251063f
c21 28 VSS 9.05081e-20
c22 29 VSS 0.00297924f
c23 30 VSS 0.014487f
r1 90 89 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r2 88 89 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r3 18 88 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3760 $Y=0.2295 $X2=0.3880 $Y2=0.2295
r4 19 18 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2295 $X2=0.3760 $Y2=0.2295
r5 84 85 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r6 86 84 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.1890 $X2=0.3635 $Y2=0.1890
r7 18 85 0.185185 $w=5.4e-08 $l=1e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r8 81 80 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r9 79 80 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4420 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r10 8 79 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4300 $Y=0.0405 $X2=0.4420 $Y2=0.0405
r11 17 8 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0405 $X2=0.4300 $Y2=0.0405
r12 16 8 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0810 $X2=0.4300 $Y2=0.0810
r13 77 16 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0810 $X2=0.4175 $Y2=0.0810
r14 73 18 15.0298 $w=2.02e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.3780 $Y=0.2045 $X2=0.3780 $Y2=0.1790
r15 7 65 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2295
+ $X2=0.3740 $Y2=0.2340
r16 7 73 14.7351 $w=2.02e-08 $l=2.5e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.3780 $Y=0.2295 $X2=0.3780 $Y2=0.2045
r17 3 59 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7830 $Y=0.1360
+ $X2=0.7830 $Y2=0.1445
r18 15 3 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=0.7830
+ $Y=0.1350 $X2=0.7830 $Y2=0.1360
r19 2 57 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7290 $Y=0.1360
+ $X2=0.7290 $Y2=0.1445
r20 14 2 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=0.7290
+ $Y=0.1350 $X2=0.7290 $Y2=0.1360
r21 8 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0405
+ $X2=0.4320 $Y2=0.0360
r22 62 63 1.98211 $w=1.3e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3830
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r23 62 65 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3830
+ $Y=0.2340 $X2=0.3740 $Y2=0.2340
r24 61 63 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r25 20 29 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4320 $Y=0.2340 $X2=0.4590 $Y2=0.2340
r26 20 61 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4050 $Y2=0.2340
r27 26 59 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1085 $X2=0.7830 $Y2=0.1445
r28 25 57 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1085 $X2=0.7290 $Y2=0.1445
r29 21 27 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4320 $Y=0.0360 $X2=0.4590 $Y2=0.0360
r30 29 50 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4590 $Y2=0.2160
r31 55 59 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.7830 $Y=0.1530
+ $X2=0.7830 $Y2=0.1445
r32 54 55 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.7560
+ $Y=0.1530 $X2=0.7830 $Y2=0.1530
r33 53 54 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1530 $X2=0.7560 $Y2=0.1530
r34 53 57 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.7290 $Y=0.1530
+ $X2=0.7290 $Y2=0.1445
r35 52 53 24.6015 $w=1.3e-08 $l=1.055e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.6235 $Y=0.1530 $X2=0.7290 $Y2=0.1530
r36 51 52 29.3819 $w=1.3e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.4975
+ $Y=0.1530 $X2=0.6235 $Y2=0.1530
r37 30 51 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M2 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1530 $X2=0.4975 $Y2=0.1530
r38 30 45 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4590 $Y=0.1530
+ $X2=0.4590 $Y2=0.1530
r39 27 44 6.39593 $w=1.55565e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4590 $Y2=0.0705
r40 49 50 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1980 $X2=0.4590 $Y2=0.2160
r41 48 49 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1800 $X2=0.4590 $Y2=0.1980
r42 47 48 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1675 $X2=0.4590 $Y2=0.1800
r43 46 47 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1630 $X2=0.4590 $Y2=0.1675
r44 45 46 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1530 $X2=0.4590 $Y2=0.1630
r45 23 45 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1415 $X2=0.4590 $Y2=0.1530
r46 23 28 1.50137 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1415 $X2=0.4590 $Y2=0.1300
r47 43 44 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1010 $X2=0.4590 $Y2=0.0705
r48 22 28 2.66732 $w=1.57273e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1135 $X2=0.4590 $Y2=0.1300
r49 22 43 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1135 $X2=0.4590 $Y2=0.1010
r50 28 41 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1300 $X2=0.4860 $Y2=0.1300
r51 40 41 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1300 $X2=0.4860 $Y2=0.1300
r52 24 38 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1300 $X2=0.5670 $Y2=0.1300
r53 24 40 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1300 $X2=0.5130 $Y2=0.1300
r54 37 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1330
+ $X2=0.5670 $Y2=0.1300
r55 1 35 0.590723 $w=1.53e-08 $l=6e-09 $layer=LIG $thickness=4.8e-08 $X=0.5670
+ $Y=0.1240 $X2=0.5670 $Y2=0.1300
r56 1 36 1.77217 $w=1.53e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08 $X=0.5670
+ $Y=0.1240 $X2=0.5670 $Y2=0.1210
r57 35 36 1.18145 $w=1.53e-08 $l=9e-09 $layer=LIG $thickness=4.8e-08 $X=0.5670
+ $Y=0.1300 $X2=0.5670 $Y2=0.1210
r58 35 37 4.72579 $w=1.53e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08 $X=0.5670
+ $Y=0.1300 $X2=0.5670 $Y2=0.1330
r59 13 35 0.314665 $w=2.27e-07 $l=5e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5670 $Y=0.1350 $X2=0.5670 $Y2=0.1300
.ends


*
.SUBCKT DHLx2_ASAP7_75t_R VSS VDD CLK D Q
*
* VSS VSS
* VDD VDD
* CLK CLK
* D D
* Q Q
*
*

MM0 N_MM0_d N_MM0_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2 N_MM2_d N_MM13_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM10_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM6 N_MM6_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM24 N_MM24_d N_MM25_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@2 N_MM24@2_d N_MM25@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM12 N_MM12_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM13 N_MM13_d N_MM13_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM25 N_MM25_d N_MM25_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@2 N_MM25@2_d N_MM25@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "DHLx2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "DHLx2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_DHLx2_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_DHLx2_ASAP7_75t_R%noxref_19
cc_1 N_noxref_19_1 N_MM3_g 0.00136823f
cc_2 N_noxref_19_1 N_CLKB_11 0.000754183f
cc_3 N_noxref_19_1 N_noxref_16_1 0.000465319f
cc_4 N_noxref_19_1 N_noxref_17_1 0.00769631f
cc_5 N_noxref_19_1 N_noxref_18_1 0.0012342f
x_PM_DHLx2_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_DHLx2_ASAP7_75t_R%noxref_18
cc_6 N_noxref_18_1 N_MM3_g 0.0013607f
cc_7 N_noxref_18_1 N_CLKB_10 0.000797943f
cc_8 N_noxref_18_1 N_noxref_16_1 0.00769877f
cc_9 N_noxref_18_1 N_noxref_17_1 0.000464978f
x_PM_DHLx2_ASAP7_75t_R%PU1 VSS N_MM3_d N_MM1_s N_PU1_1 PM_DHLx2_ASAP7_75t_R%PU1
cc_10 N_PU1_1 N_MM1_g 0.0170796f
cc_11 N_PU1_1 N_MM3_g 0.0170329f
x_PM_DHLx2_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_DHLx2_ASAP7_75t_R%noxref_15
cc_12 N_noxref_15_1 N_MM0_g 0.00367764f
cc_13 N_noxref_15_1 N_CLKN_29 5.45631e-20
cc_14 N_noxref_15_1 N_CLKN_20 8.02432e-20
cc_15 N_noxref_15_1 N_CLKN_28 8.9607e-20
cc_16 N_noxref_15_1 N_CLKN_19 0.000271574f
cc_17 N_noxref_15_1 N_CLKN_7 0.000435397f
cc_18 N_noxref_15_1 N_CLKN_18 0.0277736f
cc_19 N_noxref_15_1 N_noxref_14_1 0.0020445f
x_PM_DHLx2_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_DHLx2_ASAP7_75t_R%noxref_17
cc_20 N_noxref_17_1 N_CLKN_1 0.000395083f
cc_21 N_noxref_17_1 N_MM13_g 0.00366263f
cc_22 N_noxref_17_1 N_CLKB_11 0.0274274f
cc_23 N_noxref_17_1 N_noxref_16_1 0.00141536f
x_PM_DHLx2_ASAP7_75t_R%CLK VSS CLK N_MM0_g N_CLK_8 N_CLK_6 N_CLK_1 N_CLK_4
+ N_CLK_7 N_CLK_5 PM_DHLx2_ASAP7_75t_R%CLK
x_PM_DHLx2_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_DHLx2_ASAP7_75t_R%noxref_16
cc_24 N_noxref_16_1 N_CLKN_1 0.00039096f
cc_25 N_noxref_16_1 N_MM13_g 0.00357605f
cc_26 N_noxref_16_1 N_CLKB_10 0.0274872f
x_PM_DHLx2_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_DHLx2_ASAP7_75t_R%noxref_14
cc_27 N_noxref_14_1 N_MM0_g 0.00370865f
cc_28 N_noxref_14_1 N_CLKN_6 0.00048495f
cc_29 N_noxref_14_1 N_CLKN_27 5.82693e-20
cc_30 N_noxref_14_1 N_CLKN_19 0.000382796f
cc_31 N_noxref_14_1 N_CLKN_17 0.0276659f
x_PM_DHLx2_ASAP7_75t_R%D VSS D N_MM3_g N_D_4 N_D_1 N_D_5 PM_DHLx2_ASAP7_75t_R%D
cc_32 N_MM3_g N_CLKN_25 0.000314577f
cc_33 N_MM3_g N_CLKN_32 0.000573213f
cc_34 N_D_4 N_CLKN_33 0.000841934f
cc_35 N_D_1 N_CLKN_2 0.0023237f
cc_36 N_D_4 N_CLKN_25 0.00499725f
cc_37 N_MM3_g N_MM1_g 0.00518111f
x_PM_DHLx2_ASAP7_75t_R%PD3 VSS N_MM9_s N_MM8_d N_PD3_1 PM_DHLx2_ASAP7_75t_R%PD3
cc_38 N_PD3_1 N_MM9_g 0.00772819f
cc_39 N_PD3_1 N_MM11_g 0.00780608f
x_PM_DHLx2_ASAP7_75t_R%Q VSS Q N_MM24_d N_MM24@2_d N_MM25_d N_MM25@2_d N_Q_7
+ N_Q_9 N_Q_1 N_Q_10 N_Q_8 N_Q_2 N_Q_11 PM_DHLx2_ASAP7_75t_R%Q
cc_40 N_Q_7 N_MH_26 0.000884556f
cc_41 N_Q_7 N_MH_2 0.000493251f
cc_42 N_Q_7 N_MH_3 0.000776173f
cc_43 N_Q_9 N_MH_30 0.00123359f
cc_44 N_Q_9 N_MH_26 0.001234f
cc_45 N_Q_1 N_MH_25 0.001333f
cc_46 N_Q_10 N_MH_26 0.00139792f
cc_47 N_Q_8 N_MH_3 0.00146492f
cc_48 N_Q_8 N_MH_2 0.00159321f
cc_49 N_Q_2 N_MM25@2_g 0.00204741f
cc_50 N_Q_1 N_MM25@2_g 0.00210359f
cc_51 N_Q_11 N_MH_26 0.00535829f
cc_52 N_Q_8 N_MM25@2_g 0.0296097f
cc_53 N_Q_7 N_MM25_g 0.0368474f
cc_54 N_Q_7 N_MM25@2_g 0.0685015f
x_PM_DHLx2_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_DHLx2_ASAP7_75t_R%noxref_20
cc_55 N_noxref_20_1 N_NET088_10 0.0170016f
cc_56 N_noxref_20_1 N_MM7_g 0.00587707f
x_PM_DHLx2_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_DHLx2_ASAP7_75t_R%noxref_21
cc_57 N_noxref_21_1 N_CLKN_8 0.0028849f
cc_58 N_noxref_21_1 N_NET088_11 0.0163713f
cc_59 N_noxref_21_1 N_MM7_g 0.00529202f
cc_60 N_noxref_21_1 N_noxref_20_1 0.00147956f
x_PM_DHLx2_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_DHLx2_ASAP7_75t_R%noxref_22
cc_61 N_noxref_22_1 N_NET088_10 0.000569606f
cc_62 N_noxref_22_1 N_MM25_g 0.0016524f
cc_63 N_noxref_22_1 N_noxref_20_1 0.00775583f
cc_64 N_noxref_22_1 N_noxref_21_1 0.000452268f
x_PM_DHLx2_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_DHLx2_ASAP7_75t_R%noxref_25
cc_65 N_noxref_25_1 N_MM25@2_g 0.0015181f
cc_66 N_noxref_25_1 N_Q_8 0.000822569f
cc_67 N_noxref_25_1 N_noxref_24_1 0.00176453f
x_PM_DHLx2_ASAP7_75t_R%PD2 VSS N_MM10_s N_MM11_d N_PD2_5 N_PD2_1 N_PD2_4
+ PM_DHLx2_ASAP7_75t_R%PD2
cc_68 N_PD2_5 N_CLKN_8 0.0012587f
cc_69 N_PD2_1 N_CLKN_3 0.000885951f
cc_70 N_PD2_1 N_MM9_g 0.00219455f
cc_71 N_PD2_4 N_MM9_g 0.00714976f
cc_72 N_PD2_5 N_MM9_g 0.0240715f
cc_73 N_PD2_4 N_MM10_g 0.015035f
cc_74 N_PD2_5 N_MM11_g 0.0146095f
cc_75 N_PD2_1 N_MH_18 0.000618514f
cc_76 N_PD2_1 N_MH_20 0.000420057f
cc_77 N_PD2_1 N_MH_23 0.000432219f
cc_78 N_PD2_4 N_MH_7 0.000615363f
cc_79 N_PD2_1 N_MH_29 0.00211916f
x_PM_DHLx2_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_DHLx2_ASAP7_75t_R%noxref_23
cc_80 N_noxref_23_1 N_CLKN_8 0.00061243f
cc_81 N_noxref_23_1 N_MM25_g 0.00158717f
cc_82 N_noxref_23_1 N_noxref_20_1 0.00046976f
cc_83 N_noxref_23_1 N_noxref_21_1 0.00759211f
cc_84 N_noxref_23_1 N_noxref_22_1 0.00122968f
x_PM_DHLx2_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_DHLx2_ASAP7_75t_R%noxref_24
cc_85 N_noxref_24_1 N_MM25@2_g 0.00153744f
cc_86 N_noxref_24_1 N_Q_7 0.000822557f
x_PM_DHLx2_ASAP7_75t_R%PD1 VSS N_MM5_d N_MM4_s N_PD1_5 N_PD1_4 N_PD1_1
+ PM_DHLx2_ASAP7_75t_R%PD1
cc_87 N_PD1_5 N_CLKN_25 0.000471129f
cc_88 N_PD1_5 N_CLKN_2 0.00249638f
cc_89 N_PD1_5 N_MM1_g 0.0737346f
cc_90 N_PD1_4 N_D_1 0.000644276f
cc_91 N_PD1_4 N_D_4 0.000738512f
cc_92 N_PD1_4 N_MM3_g 0.0361099f
cc_93 N_PD1_5 N_CLKB_1 0.000659769f
cc_94 N_PD1_5 N_MM10_g 0.0347952f
cc_95 N_PD1_1 N_MH_21 0.000163055f
cc_96 N_PD1_1 N_MH_8 0.00139646f
cc_97 N_PD1_1 N_MH_16 0.00319382f
x_PM_DHLx2_ASAP7_75t_R%CLKN VSS N_MM13_g N_MM1_g N_MM9_g N_MM0_d N_MM12_d
+ N_CLKN_31 N_CLKN_24 N_CLKN_28 N_CLKN_30 N_CLKN_7 N_CLKN_6 N_CLKN_17 N_CLKN_18
+ N_CLKN_1 N_CLKN_22 N_CLKN_19 N_CLKN_23 N_CLKN_33 N_CLKN_21 N_CLKN_25
+ N_CLKN_32 N_CLKN_2 N_CLKN_8 N_CLKN_3 N_CLKN_26 N_CLKN_27 N_CLKN_29 N_CLKN_20
+ PM_DHLx2_ASAP7_75t_R%CLKN
cc_98 N_CLKN_31 N_MM0_g 9.71373e-20
cc_99 N_CLKN_24 N_MM0_g 0.000107013f
cc_100 N_CLKN_28 N_MM0_g 0.000184097f
cc_101 N_CLKN_30 N_MM0_g 0.000187475f
cc_102 N_CLKN_7 N_MM0_g 0.00107419f
cc_103 N_CLKN_6 N_MM0_g 0.00115113f
cc_104 N_CLKN_17 N_MM0_g 0.0112216f
cc_105 N_CLKN_18 N_MM0_g 0.0113259f
cc_106 N_CLKN_1 N_CLK_8 0.000441107f
cc_107 N_CLKN_22 N_CLK_6 0.000655904f
cc_108 N_CLKN_1 N_CLK_1 0.00331106f
cc_109 N_CLKN_19 N_CLK_4 0.00106325f
cc_110 N_CLKN_23 N_CLK_8 0.00120365f
cc_111 N_CLKN_23 N_CLK_7 0.00139663f
cc_112 N_CLKN_30 N_CLK_8 0.00151884f
cc_113 N_CLKN_33 N_CLK_6 0.0017293f
cc_114 N_CLKN_21 N_CLK_5 0.001733f
cc_115 N_CLKN_30 N_CLK_6 0.00235877f
cc_116 N_CLKN_28 N_CLK_8 0.0029115f
cc_117 N_CLKN_19 N_CLK_7 0.00295223f
cc_118 N_MM13_g N_MM0_g 0.0351254f
x_PM_DHLx2_ASAP7_75t_R%NET088 VSS N_MM11_g N_MM6_d N_MM7_d N_NET088_11
+ N_NET088_16 N_NET088_1 N_NET088_4 N_NET088_14 N_NET088_3 N_NET088_13
+ N_NET088_15 N_NET088_10 N_NET088_12 PM_DHLx2_ASAP7_75t_R%NET088
cc_119 N_MM11_g N_CLKN_8 0.00513228f
cc_120 N_MM11_g N_CLKN_3 0.000148702f
cc_121 N_MM11_g N_CLKN_33 0.000207036f
cc_122 N_MM11_g N_CLKN_26 0.000291947f
cc_123 N_NET088_11 N_CLKN_8 0.000379755f
cc_124 N_NET088_16 N_CLKN_8 0.000406877f
cc_125 N_NET088_1 N_MM9_g 0.00042377f
cc_126 N_NET088_4 N_CLKN_8 0.000892611f
cc_127 N_NET088_14 N_CLKN_8 0.00135202f
cc_128 N_MM11_g N_MM9_g 0.0144008f
x_PM_DHLx2_ASAP7_75t_R%CLKB VSS N_MM10_g N_MM2_d N_MM13_d N_CLKB_3 N_CLKB_4
+ N_CLKB_13 N_CLKB_12 N_CLKB_10 N_CLKB_11 N_CLKB_18 N_CLKB_15 N_CLKB_14
+ N_CLKB_1 N_CLKB_17 N_CLKB_16 PM_DHLx2_ASAP7_75t_R%CLKB
cc_129 N_CLKB_3 N_CLK_5 0.000437879f
cc_130 N_CLKB_4 N_CLK_5 0.00019816f
cc_131 N_CLKB_13 N_CLK_6 0.00106614f
cc_132 N_CLKB_12 N_CLK_5 0.00272143f
cc_133 N_CLKB_10 N_CLKN_19 5.89059e-20
cc_134 N_CLKB_10 N_CLKN_8 0.000115256f
cc_135 N_CLKB_10 N_CLKN_30 0.000221545f
cc_136 N_CLKB_4 N_CLKN_30 0.000283373f
cc_137 N_CLKB_13 N_CLKN_30 0.00474673f
cc_138 N_CLKB_11 N_MM13_g 0.0111457f
cc_139 N_CLKB_18 N_CLKN_25 0.000395204f
cc_140 N_CLKB_4 N_CLKN_1 0.000415101f
cc_141 N_CLKB_12 N_CLKN_31 0.000487526f
cc_142 N_CLKB_15 N_CLKN_32 0.000492957f
cc_143 N_CLKB_14 N_CLKN_23 0.000601159f
cc_144 N_CLKB_15 N_CLKN_33 0.000665257f
cc_145 N_MM10_g N_CLKN_3 0.000675128f
cc_146 N_CLKB_3 N_MM13_g 0.00074301f
cc_147 N_CLKB_11 N_CLKN_1 0.000901256f
cc_148 N_CLKB_1 N_CLKN_2 0.00226448f
cc_149 N_CLKB_14 N_CLKN_33 0.000938226f
cc_150 N_CLKB_4 N_MM13_g 0.00111127f
cc_151 N_CLKB_14 N_CLKN_24 0.0011563f
cc_152 N_MM10_g N_MM1_g 0.00162675f
cc_153 N_CLKB_15 N_CLKN_25 0.00354617f
cc_154 N_CLKB_14 N_CLKN_31 0.00377879f
cc_155 N_MM10_g N_MM9_g 0.00908419f
cc_156 N_CLKB_18 N_CLKN_33 0.0194855f
cc_157 N_CLKB_10 N_MM13_g 0.0389364f
cc_158 N_CLKB_17 N_D_4 0.000307404f
cc_159 N_CLKB_16 N_D_5 0.000948602f
cc_160 N_CLKB_18 N_D_4 0.00106517f
cc_161 N_CLKB_14 N_D_4 0.00851671f
x_PM_DHLx2_ASAP7_75t_R%MH VSS N_MM7_g N_MM25_g N_MM25@2_g N_MM4_d N_MM9_d
+ N_MM1_d N_MM10_d N_MH_16 N_MH_20 N_MH_19 N_MH_17 N_MH_22 N_MH_7 N_MH_18
+ N_MH_29 N_MH_23 N_MH_1 N_MH_30 N_MH_24 N_MH_8 N_MH_21 N_MH_28 N_MH_2 N_MH_25
+ N_MH_27 N_MH_26 N_MH_3 PM_DHLx2_ASAP7_75t_R%MH
cc_162 N_MH_16 N_CLKN_26 0.000124991f
cc_163 N_MH_20 N_CLKN_25 0.000132722f
cc_164 N_MH_19 N_MM1_g 0.000151732f
cc_165 N_MH_17 N_MM9_g 0.000170254f
cc_166 N_MH_22 N_CLKN_26 0.000243602f
cc_167 N_MH_7 N_CLKN_2 0.000250516f
cc_168 N_MH_18 N_MM1_g 0.0346117f
cc_169 N_MH_7 N_CLKN_32 0.000312376f
cc_170 N_MH_29 N_CLKN_26 0.000411728f
cc_171 N_MH_23 N_CLKN_33 0.000468675f
cc_172 N_MH_7 N_CLKN_25 0.000516723f
cc_173 N_MH_1 N_CLKN_8 0.00175356f
cc_174 N_MH_30 N_CLKN_26 0.000650185f
cc_175 N_MH_24 N_CLKN_8 0.000651709f
cc_176 N_MH_8 N_MM9_g 0.000660894f
cc_177 N_MH_18 N_CLKN_2 0.000774744f
cc_178 N_MH_23 N_CLKN_3 0.000929711f
cc_179 N_MH_7 N_MM1_g 0.00194946f
cc_180 N_MH_24 N_CLKN_26 0.00205617f
cc_181 N_MH_20 N_CLKN_32 0.00364433f
cc_182 N_MH_30 N_CLKN_33 0.00457893f
cc_183 N_MH_23 N_CLKN_26 0.00460911f
cc_184 N_MH_20 N_CLKN_33 0.00570508f
cc_185 N_MM7_g N_CLKN_8 0.00630582f
cc_186 N_MH_16 N_MM9_g 0.0370448f
cc_187 N_MH_17 N_MM10_g 0.000138687f
cc_188 N_MH_19 N_MM10_g 0.000177764f
cc_189 N_MH_21 N_CLKB_15 0.000245663f
cc_190 N_MH_20 N_CLKB_15 0.000297537f
cc_191 N_MH_18 N_MM10_g 0.0167631f
cc_192 N_MH_30 N_CLKB_18 0.000649273f
cc_193 N_MH_23 N_CLKB_15 0.00176797f
cc_194 N_MH_22 N_CLKB_15 0.000852604f
cc_195 N_MH_20 N_CLKB_18 0.000884406f
cc_196 N_MH_8 N_CLKB_1 0.000896545f
cc_197 N_MH_8 N_MM10_g 0.0011185f
cc_198 N_MH_7 N_MM10_g 0.00118512f
cc_199 N_MH_16 N_CLKB_1 0.00170397f
cc_200 N_MH_28 N_CLKB_15 0.00285843f
cc_201 N_MH_16 N_MM10_g 0.0538222f
cc_202 N_MH_2 N_MM11_g 0.000141072f
cc_203 N_MH_21 N_MM11_g 7.10339e-20
cc_204 N_MH_25 N_MM11_g 8.03079e-20
cc_205 N_MH_16 N_MM11_g 0.000168632f
cc_206 N_MH_24 N_MM11_g 0.000173219f
cc_207 N_MM7_g N_NET088_11 0.00678056f
cc_208 N_MM7_g N_NET088_3 0.000363693f
cc_209 N_MH_30 N_NET088_16 0.000434718f
cc_210 N_MH_8 N_NET088_1 0.000438812f
cc_211 N_MH_25 N_NET088_14 0.000454057f
cc_212 N_MH_24 N_NET088_13 0.000614094f
cc_213 N_MH_1 N_NET088_14 0.000798657f
cc_214 N_MH_27 N_NET088_15 0.000912245f
cc_215 N_MH_24 N_NET088_1 0.000923139f
cc_216 N_MH_1 N_MM11_g 0.000927203f
cc_217 N_MM7_g N_NET088_1 0.00108474f
cc_218 N_MM7_g N_NET088_10 0.00660824f
cc_219 N_MH_30 N_NET088_14 0.0025869f
cc_220 N_MH_24 N_NET088_12 0.00301942f
cc_221 N_MH_22 N_NET088_12 0.00362099f
cc_222 N_MH_24 N_NET088_14 0.00404733f
cc_223 N_MM7_g N_MM11_g 0.0291006f
*END of DHLx2_ASAP7_75t_R.pxi
.ENDS
** Design:	DHLx3_ASAP7_75t_R
* Created:	"Fri Aug 17 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "DHLx3_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "DHLx3_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_DHLx3_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.0418477f
.ends

.subckt PM_DHLx3_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.0419127f
.ends

.subckt PM_DHLx3_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00432978f
.ends

.subckt PM_DHLx3_ASAP7_75t_R%PD3 VSS 2 4 1
c1 1 VSS 0.000878943f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0405 $X2=0.4905 $Y2=0.0405
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0405 $X2=0.4735 $Y2=0.0405
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4735 $Y=0.0405 $X2=0.4905 $Y2=0.0405
.ends

.subckt PM_DHLx3_ASAP7_75t_R%CLK VSS 11 3 8 6 1 4 7 5
c1 1 VSS 0.00253523f
c2 3 VSS 0.0596883f
c3 4 VSS 0.000762511f
c4 5 VSS 0.00428688f
c5 6 VSS 0.00416706f
c6 7 VSS 0.00189244f
c7 8 VSS 0.00164398f
r1 6 17 1.35805 $w=2.83333e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.1935 $X2=0.1080 $Y2=0.1710
r2 5 15 4.50612 $w=2.06667e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0630 $X2=0.1080 $Y2=0.0990
r3 16 17 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.1710 $X2=0.1080 $Y2=0.1710
r4 8 13 1.35805 $w=2.83333e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1710 $X2=0.0810 $Y2=0.1485
r5 8 16 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1710 $X2=0.0945 $Y2=0.1710
r6 14 15 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.0990 $X2=0.1080 $Y2=0.0990
r7 7 10 0.483592 $w=3.42308e-08 $l=1.87e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0990 $X2=0.0810 $Y2=0.1177
r8 7 14 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0990 $X2=0.0945 $Y2=0.0990
r9 11 12 0.874462 $w=1.3e-08 $l=3.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1227
r10 11 10 0.291487 $w=1.3e-08 $l=1.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1177
r11 4 12 2.85657 $w=1.3e-08 $l=1.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1227
r12 4 13 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1485
r13 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r14 1 4 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_DHLx3_ASAP7_75t_R%PU1 VSS 2 4 1
c1 1 VSS 0.000967541f
r1 4 3 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3365 $Y2=0.2025
r2 2 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3195 $Y2=0.2025
r3 1 3 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3195 $Y=0.2025 $X2=0.3365 $Y2=0.2025
.ends

.subckt PM_DHLx3_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00423907f
.ends

.subckt PM_DHLx3_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.00475267f
.ends

.subckt PM_DHLx3_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.00469298f
.ends

.subckt PM_DHLx3_ASAP7_75t_R%D VSS 9 3 4 1 5
c1 1 VSS 0.00711602f
c2 3 VSS 0.0838904f
c3 4 VSS 0.00909584f
c4 5 VSS 0.00704778f
r1 10 11 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1215 $X2=0.2970 $Y2=0.1350
r2 9 10 1.16595 $w=1.3e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1165 $X2=0.2970 $Y2=0.1215
r3 9 8 1.28254 $w=1.3e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1165 $X2=0.2970 $Y2=0.1110
r4 4 8 8.27824 $w=1.3e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0755 $X2=0.2970 $Y2=0.1110
r5 4 5 8.03069 $w=1.41392e-08 $l=3.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0755 $X2=0.2970 $Y2=0.0360
r6 3 1 6.51726 $w=1.18568e-07 $l=5e-10 $layer=LIG $thickness=5.19024e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2970 $Y2=0.1345
r7 1 11 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1345
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_DHLx3_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.0034898f
.ends

.subckt PM_DHLx3_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.00390159f
.ends

.subckt PM_DHLx3_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.00534346f
.ends

.subckt PM_DHLx3_ASAP7_75t_R%NET29 VSS 9 35 41 4 11 16 1 14 3 13 15 10 12 17
c1 1 VSS 0.0028932f
c2 3 VSS 0.00568573f
c3 4 VSS 0.00641745f
c4 9 VSS 0.0375042f
c5 10 VSS 0.00320676f
c6 11 VSS 0.00339735f
c7 12 VSS 0.00128775f
c8 13 VSS 0.0083537f
c9 14 VSS 0.0028093f
c10 15 VSS 0.00342499f
c11 16 VSS 0.00632305f
c12 17 VSS 0.0024621f
r1 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2295 $X2=0.5920 $Y2=0.2295
r2 41 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.2295 $X2=0.5795 $Y2=0.2295
r3 4 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2295
+ $X2=0.5940 $Y2=0.2340
r4 37 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.2340 $X2=0.6075 $Y2=0.2340
r5 16 33 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.2340 $X2=0.6210 $Y2=0.2160
r6 16 38 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.2340 $X2=0.6075 $Y2=0.2340
r7 10 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.0405 $X2=0.5920 $Y2=0.0405
r8 35 10 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0405 $X2=0.5795 $Y2=0.0405
r9 32 33 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1870 $X2=0.6210 $Y2=0.2160
r10 31 32 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1655 $X2=0.6210 $Y2=0.1870
r11 30 31 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1515 $X2=0.6210 $Y2=0.1655
r12 29 30 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1300 $X2=0.6210 $Y2=0.1515
r13 28 29 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1085 $X2=0.6210 $Y2=0.1300
r14 27 28 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0930 $X2=0.6210 $Y2=0.1085
r15 14 17 5.69636 $w=1.58e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.0675 $X2=0.6210 $Y2=0.0360
r16 14 27 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0675 $X2=0.6210 $Y2=0.0930
r17 3 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0405
+ $X2=0.5940 $Y2=0.0360
r18 17 26 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.0360 $X2=0.6075 $Y2=0.0360
r19 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0360 $X2=0.6075 $Y2=0.0360
r20 24 25 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5830
+ $Y=0.0360 $X2=0.5940 $Y2=0.0360
r21 13 15 7.32869 $w=1.41688e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5515 $Y=0.0360 $X2=0.5130 $Y2=0.0360
r22 13 24 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5515
+ $Y=0.0360 $X2=0.5830 $Y2=0.0360
r23 12 22 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0590 $X2=0.5130 $Y2=0.0820
r24 12 15 3.71425 $w=1.68348e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.0590 $X2=0.5130 $Y2=0.0360
r25 1 19 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.5130
+ $Y=0.0820 $X2=0.5130 $Y2=0.0820
r26 1 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.0820
+ $X2=0.5130 $Y2=0.0820
r27 9 19 0.314665 $w=2.27e-07 $l=5.3e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5130 $Y2=0.0820
.ends

.subckt PM_DHLx3_ASAP7_75t_R%PD2 VSS 7 13 4 5 1
c1 1 VSS 0.00756023f
c2 4 VSS 0.00184274f
c3 5 VSS 0.00233271f
r1 13 12 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r2 5 12 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4880 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r3 10 5 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4725
+ $Y=0.2295 $X2=0.4860 $Y2=0.2295
r4 9 10 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4590
+ $Y=0.2295 $X2=0.4725 $Y2=0.2295
r5 8 9 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4455
+ $Y=0.2295 $X2=0.4590 $Y2=0.2295
r6 1 8 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4320
+ $Y=0.2295 $X2=0.4455 $Y2=0.2295
r7 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2295 $X2=0.4300 $Y2=0.2295
r8 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2295 $X2=0.4175 $Y2=0.2295
.ends

.subckt PM_DHLx3_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.042337f
.ends

.subckt PM_DHLx3_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.0423286f
.ends

.subckt PM_DHLx3_ASAP7_75t_R%PD1 VSS 7 10 4 5 1
c1 1 VSS 0.0096015f
c2 4 VSS 0.00314457f
c3 5 VSS 0.00187694f
r1 10 9 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r2 8 9 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r3 5 8 0.123457 $w=8.1e-08 $l=1e-08 $layer=N_src_drn $thickness=1e-09 $X=0.3780
+ $Y=0.0675 $X2=0.3880 $Y2=0.0675
r4 4 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3220 $Y2=0.0675
r5 7 4 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r6 1 5 1e-05
.ends

.subckt PM_DHLx3_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.00535381f
.ends

.subckt PM_DHLx3_ASAP7_75t_R%Q VSS 42 23 39 40 62 63 65 1 18 17 2 14 3 15 13 19
+ 4 16
c1 1 VSS 0.00820532f
c2 2 VSS 0.00832217f
c3 3 VSS 0.00994934f
c4 4 VSS 0.00980191f
c5 13 VSS 0.00341783f
c6 14 VSS 0.00448051f
c7 15 VSS 0.00394137f
c8 16 VSS 0.00446565f
c9 17 VSS 0.0182852f
c10 18 VSS 0.0173352f
c11 19 VSS 0.00667036f
c12 20 VSS 0.00313114f
c13 21 VSS 0.00330069f
r1 65 64 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.2025 $X2=0.7165 $Y2=0.2025
r2 15 64 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7040 $Y=0.2025 $X2=0.7165 $Y2=0.2025
r3 63 61 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8270 $Y=0.2025 $X2=0.8245 $Y2=0.2025
r4 4 61 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8100 $Y=0.2025 $X2=0.8245 $Y2=0.2025
r5 16 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.2025 $X2=0.8100 $Y2=0.2025
r6 62 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.2025 $X2=0.7955 $Y2=0.2025
r7 2 53 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7020 $Y=0.2295
+ $X2=0.7020 $Y2=0.2340
r8 4 47 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8100 $Y=0.2025
+ $X2=0.8100 $Y2=0.2340
r9 53 54 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.2340 $X2=0.7155 $Y2=0.2340
r10 51 54 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.2340 $X2=0.7155 $Y2=0.2340
r11 50 51 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.2340 $X2=0.7290 $Y2=0.2340
r12 49 50 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.2340 $X2=0.7560 $Y2=0.2340
r13 47 48 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.2340 $X2=0.8235 $Y2=0.2340
r14 46 47 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7965
+ $Y=0.2340 $X2=0.8100 $Y2=0.2340
r15 46 49 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7965
+ $Y=0.2340 $X2=0.7830 $Y2=0.2340
r16 45 48 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.2340 $X2=0.8235 $Y2=0.2340
r17 18 21 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8640 $Y=0.2340 $X2=0.8910 $Y2=0.2340
r18 18 45 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.2340 $X2=0.8370 $Y2=0.2340
r19 21 44 7.2121 $w=1.53211e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8910 $Y=0.2340 $X2=0.8910 $Y2=0.1960
r20 43 44 8.33653 $w=1.3e-08 $l=3.58e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1602 $X2=0.8910 $Y2=0.1960
r21 42 43 1.69063 $w=1.3e-08 $l=7.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1530 $X2=0.8910 $Y2=0.1602
r22 42 41 7.40378 $w=1.3e-08 $l=3.18e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1530 $X2=0.8910 $Y2=0.1212
r23 19 20 5.69636 $w=1.58e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8910 $Y=0.0675 $X2=0.8910 $Y2=0.0360
r24 19 41 12.5339 $w=1.3e-08 $l=5.37e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.0675 $X2=0.8910 $Y2=0.1212
r25 40 38 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8270 $Y=0.0675 $X2=0.8245 $Y2=0.0675
r26 3 38 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8100 $Y=0.0675 $X2=0.8245 $Y2=0.0675
r27 14 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.0675 $X2=0.8100 $Y2=0.0675
r28 39 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.0675 $X2=0.7955 $Y2=0.0675
r29 20 36 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8910 $Y=0.0360 $X2=0.8640 $Y2=0.0360
r30 3 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8100 $Y=0.0675
+ $X2=0.8100 $Y2=0.0360
r31 35 36 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.0360 $X2=0.8640 $Y2=0.0360
r32 34 35 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8235
+ $Y=0.0360 $X2=0.8370 $Y2=0.0360
r33 33 34 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0360 $X2=0.8235 $Y2=0.0360
r34 32 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7965
+ $Y=0.0360 $X2=0.8100 $Y2=0.0360
r35 31 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.0360 $X2=0.7965 $Y2=0.0360
r36 30 31 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.0360 $X2=0.7830 $Y2=0.0360
r37 29 30 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.0360 $X2=0.7560 $Y2=0.0360
r38 28 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7155
+ $Y=0.0360 $X2=0.7290 $Y2=0.0360
r39 27 28 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.0360 $X2=0.7155 $Y2=0.0360
r40 17 27 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6905
+ $Y=0.0360 $X2=0.7020 $Y2=0.0360
r41 13 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7020 $Y=0.0405
+ $X2=0.7020 $Y2=0.0360
r42 1 13 12.9669 $w=2.02e-08 $l=2.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7020 $Y=0.0625 $X2=0.7020 $Y2=0.0405
r43 23 22 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.0675 $X2=0.7165 $Y2=0.0675
r44 13 22 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7040 $Y=0.0675 $X2=0.7165 $Y2=0.0675
r45 2 15 1e-05
.ends

.subckt PM_DHLx3_ASAP7_75t_R%MH VSS 15 16 17 18 88 92 98 102 23 32 22 20 9 25
+ 21 33 1 26 10 34 27 19 24 28 2 31 30 29 3 4
c1 1 VSS 0.00034616f
c2 2 VSS 0.00415614f
c3 3 VSS 0.00382455f
c4 4 VSS 0.00387055f
c5 9 VSS 0.00632495f
c6 10 VSS 0.00511036f
c7 15 VSS 0.0368895f
c8 16 VSS 0.0800705f
c9 17 VSS 0.0801427f
c10 18 VSS 0.0804318f
c11 19 VSS 0.00521728f
c12 20 VSS 0.00143536f
c13 21 VSS 0.00556032f
c14 22 VSS 0.0014312f
c15 23 VSS 0.00837554f
c16 24 VSS 0.00410433f
c17 25 VSS 0.00141777f
c18 26 VSS 0.000757319f
c19 27 VSS 0.000517962f
c20 28 VSS 0.00247731f
c21 29 VSS 0.00222214f
c22 30 VSS 0.00291916f
c23 31 VSS 0.00332151f
c24 32 VSS 7.84211e-20
c25 33 VSS 0.00250514f
c26 34 VSS 0.0195804f
r1 102 101 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r2 100 101 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r3 21 100 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3760 $Y=0.2295 $X2=0.3880 $Y2=0.2295
r4 22 21 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2295 $X2=0.3760 $Y2=0.2295
r5 96 97 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r6 98 96 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.1890 $X2=0.3635 $Y2=0.1890
r7 21 97 0.185185 $w=5.4e-08 $l=1e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r8 92 91 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r9 90 91 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4420 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r10 10 90 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4300 $Y=0.0405 $X2=0.4420 $Y2=0.0405
r11 20 10 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0405 $X2=0.4300 $Y2=0.0405
r12 19 10 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0810 $X2=0.4300 $Y2=0.0810
r13 88 19 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0810 $X2=0.4175 $Y2=0.0810
r14 84 21 15.0298 $w=2.02e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.3780 $Y=0.2045 $X2=0.3780 $Y2=0.1790
r15 9 74 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2295
+ $X2=0.3740 $Y2=0.2340
r16 9 84 14.7351 $w=2.02e-08 $l=2.5e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.3780 $Y=0.2295 $X2=0.3780 $Y2=0.2045
r17 4 68 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8370 $Y=0.1360
+ $X2=0.8370 $Y2=0.1445
r18 18 4 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=0.8370
+ $Y=0.1350 $X2=0.8370 $Y2=0.1360
r19 3 66 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7830 $Y=0.1360
+ $X2=0.7830 $Y2=0.1445
r20 17 3 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=0.7830
+ $Y=0.1350 $X2=0.7830 $Y2=0.1360
r21 2 64 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7290 $Y=0.1360
+ $X2=0.7290 $Y2=0.1445
r22 16 2 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=0.7290
+ $Y=0.1350 $X2=0.7290 $Y2=0.1360
r23 10 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0405
+ $X2=0.4320 $Y2=0.0360
r24 71 72 1.98211 $w=1.3e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3830
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r25 71 74 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3830
+ $Y=0.2340 $X2=0.3740 $Y2=0.2340
r26 70 72 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r27 23 33 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4320 $Y=0.2340 $X2=0.4590 $Y2=0.2340
r28 23 70 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4050 $Y2=0.2340
r29 30 68 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1085 $X2=0.8370 $Y2=0.1445
r30 29 66 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1085 $X2=0.7830 $Y2=0.1445
r31 28 64 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1085 $X2=0.7290 $Y2=0.1445
r32 24 31 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4320 $Y=0.0360 $X2=0.4590 $Y2=0.0360
r33 33 55 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4590 $Y2=0.2160
r34 62 68 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.8370 $Y=0.1530
+ $X2=0.8370 $Y2=0.1445
r35 61 62 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.8100
+ $Y=0.1530 $X2=0.8370 $Y2=0.1530
r36 60 61 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1530 $X2=0.8100 $Y2=0.1530
r37 60 66 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.7830 $Y=0.1530
+ $X2=0.7830 $Y2=0.1445
r38 59 60 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.7560
+ $Y=0.1530 $X2=0.7830 $Y2=0.1530
r39 58 59 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1530 $X2=0.7560 $Y2=0.1530
r40 58 64 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.7290 $Y=0.1530
+ $X2=0.7290 $Y2=0.1445
r41 57 58 24.6015 $w=1.3e-08 $l=1.055e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.6235 $Y=0.1530 $X2=0.7290 $Y2=0.1530
r42 56 57 29.3819 $w=1.3e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.4975
+ $Y=0.1530 $X2=0.6235 $Y2=0.1530
r43 34 56 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M2 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1530 $X2=0.4975 $Y2=0.1530
r44 34 50 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4590 $Y=0.1530
+ $X2=0.4590 $Y2=0.1530
r45 31 49 6.39593 $w=1.55565e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4590 $Y2=0.0705
r46 54 55 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1980 $X2=0.4590 $Y2=0.2160
r47 53 54 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1800 $X2=0.4590 $Y2=0.1980
r48 52 53 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1675 $X2=0.4590 $Y2=0.1800
r49 51 52 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1630 $X2=0.4590 $Y2=0.1675
r50 50 51 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1530 $X2=0.4590 $Y2=0.1630
r51 26 50 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1415 $X2=0.4590 $Y2=0.1530
r52 26 32 1.50137 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1415 $X2=0.4590 $Y2=0.1300
r53 48 49 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1010 $X2=0.4590 $Y2=0.0705
r54 25 32 2.66732 $w=1.57273e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1135 $X2=0.4590 $Y2=0.1300
r55 25 48 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1135 $X2=0.4590 $Y2=0.1010
r56 32 46 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1300 $X2=0.4860 $Y2=0.1300
r57 45 46 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1300 $X2=0.4860 $Y2=0.1300
r58 27 43 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1300 $X2=0.5670 $Y2=0.1300
r59 27 45 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1300 $X2=0.5130 $Y2=0.1300
r60 42 43 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1330
+ $X2=0.5670 $Y2=0.1300
r61 1 40 0.590723 $w=1.53e-08 $l=6e-09 $layer=LIG $thickness=4.8e-08 $X=0.5670
+ $Y=0.1240 $X2=0.5670 $Y2=0.1300
r62 1 41 1.77217 $w=1.53e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08 $X=0.5670
+ $Y=0.1240 $X2=0.5670 $Y2=0.1210
r63 40 41 1.18145 $w=1.53e-08 $l=9e-09 $layer=LIG $thickness=4.8e-08 $X=0.5670
+ $Y=0.1300 $X2=0.5670 $Y2=0.1210
r64 40 42 4.72579 $w=1.53e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08 $X=0.5670
+ $Y=0.1300 $X2=0.5670 $Y2=0.1330
r65 15 40 0.314665 $w=2.27e-07 $l=5e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5670 $Y=0.1350 $X2=0.5670 $Y2=0.1300
.ends

.subckt PM_DHLx3_ASAP7_75t_R%CLKN VSS 14 15 16 99 101 24 31 28 30 7 6 18 17 1
+ 22 19 23 33 21 32 2 25 8 3 26 27 29 20
c1 1 VSS 0.00164427f
c2 2 VSS 0.000269886f
c3 3 VSS 0.000104638f
c4 6 VSS 0.00755633f
c5 7 VSS 0.00768933f
c6 8 VSS 0.00485057f
c7 14 VSS 0.059914f
c8 15 VSS 0.00535598f
c9 16 VSS 0.00506338f
c10 17 VSS 0.00583713f
c11 18 VSS 0.00576435f
c12 19 VSS 0.00681165f
c13 20 VSS 0.00154771f
c14 21 VSS 0.00491212f
c15 22 VSS 0.00378952f
c16 23 VSS 0.000478308f
c17 24 VSS 0.000243113f
c18 25 VSS 0.000859229f
c19 26 VSS 0.00158728f
c20 27 VSS 0.00353633f
c21 28 VSS 0.00157772f
c22 29 VSS 0.00370372f
c23 30 VSS 0.000777959f
c24 31 VSS 0.000467133f
c25 32 VSS 0.000588563f
c26 33 VSS 0.0206551f
r1 101 100 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r2 18 100 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r3 99 98 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r4 17 98 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r5 7 96 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0550 $Y2=0.2340
r6 6 93 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0550 $Y2=0.0360
r7 95 96 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.2340 $X2=0.0550 $Y2=0.2340
r8 22 95 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0460 $Y2=0.2340
r9 22 29 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0180 $Y2=0.2340
r10 92 93 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.0360 $X2=0.0550 $Y2=0.0360
r11 21 92 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0460 $Y2=0.0360
r12 21 27 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0180 $Y2=0.0360
r13 3 82 5.67512 $w=2.4e-08 $l=5e-09 $layer=LISD $thickness=4.02632e-08
+ $X=0.4590 $Y=0.1790 $X2=0.4640 $Y2=0.1790
r14 16 3 2.88446 $w=1.16273e-07 $l=4.4e-08 $layer=LIG $thickness=5.16364e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4590 $Y2=0.1790
r15 15 76 6.51726 $w=1.18568e-07 $l=5e-10 $layer=LIG $thickness=5.19024e-08
+ $X=0.3510 $Y=0.1350 $X2=0.3510 $Y2=0.1345
r16 27 75 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.0360 $X2=0.0180 $Y2=0.0630
r17 80 82 11.0623 $w=2.14976e-08 $l=2.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4845 $Y=0.1790 $X2=0.4640 $Y2=0.1790
r18 79 80 8.84105 $w=2.02e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4995 $Y=0.1790 $X2=0.4845 $Y2=0.1790
r19 8 77 6.18874 $w=2.02e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5025 $Y=0.1790 $X2=0.5130 $Y2=0.1790
r20 8 79 1.76821 $w=2.02e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.5025
+ $Y=0.1790 $X2=0.4995 $Y2=0.1790
r21 2 76 6.49795 $w=1.53e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08 $X=0.3510
+ $Y=0.1235 $X2=0.3510 $Y2=0.1345
r22 20 28 3.9134 $w=1.47857e-08 $l=2.25499e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.2115 $X2=0.0165 $Y2=0.1890
r23 20 29 3.59766 $w=1.692e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.2115 $X2=0.0180 $Y2=0.2340
r24 74 75 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0990 $X2=0.0180 $Y2=0.0630
r25 73 74 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1350 $X2=0.0180 $Y2=0.0990
r26 19 28 3.9134 $w=1.47857e-08 $l=2.25499e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1665 $X2=0.0165 $Y2=0.1890
r27 19 73 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1665 $X2=0.0180 $Y2=0.1350
r28 71 77 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5130 $Y=0.1845
+ $X2=0.5130 $Y2=0.1790
r29 26 71 3.96423 $w=1.3e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1675 $X2=0.5130 $Y2=0.1845
r30 32 65 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.1980 $X2=0.3510 $Y2=0.1845
r31 32 56 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.3510 $Y=0.1980 $X2=0.3510
+ $Y2=0.1890
r32 67 68 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1340 $X2=0.3510 $Y2=0.1570
r33 67 76 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1340
+ $X2=0.3510 $Y2=0.1345
r34 25 65 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1755 $X2=0.3510 $Y2=0.1845
r35 25 68 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1755 $X2=0.3510 $Y2=0.1570
r36 62 63 1.90199 $w=1.38333e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.0255 $Y=0.1890 $X2=0.0345 $Y2=0.1890
r37 28 62 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0165
+ $Y=0.1890 $X2=0.0255 $Y2=0.1890
r38 60 71 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.5130 $Y=0.1890
+ $X2=0.5130 $Y2=0.1845
r39 59 60 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.4770
+ $Y=0.1890 $X2=0.5130 $Y2=0.1890
r40 58 59 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M2 $thickness=3.6e-08 $X=0.4320
+ $Y=0.1890 $X2=0.4770 $Y2=0.1890
r41 57 58 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M2 $thickness=3.6e-08 $X=0.3870
+ $Y=0.1890 $X2=0.4320 $Y2=0.1890
r42 56 57 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1890 $X2=0.3870 $Y2=0.1890
r43 56 65 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.3510 $Y=0.1890 $X2=0.3510
+ $Y2=0.1845
r44 55 56 15.2739 $w=1.3e-08 $l=6.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.2855
+ $Y=0.1890 $X2=0.3510 $Y2=0.1890
r45 54 55 19.9377 $w=1.3e-08 $l=8.55e-08 $layer=M2 $thickness=3.6e-08 $X=0.2000
+ $Y=0.1890 $X2=0.2855 $Y2=0.1890
r46 53 54 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.1620
+ $Y=0.1890 $X2=0.2000 $Y2=0.1890
r47 52 53 15.0407 $w=1.3e-08 $l=6.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.0975
+ $Y=0.1890 $X2=0.1620 $Y2=0.1890
r48 51 52 15.0407 $w=1.3e-08 $l=6.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.0330
+ $Y=0.1890 $X2=0.0975 $Y2=0.1890
r49 51 63 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.0330 $Y=0.1890
+ $X2=0.0345 $Y2=0.1890
r50 33 51 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.0215
+ $Y=0.1890 $X2=0.0330 $Y2=0.1890
r51 49 50 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.1890 $X2=0.1755 $Y2=0.1890
r52 49 53 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1620 $Y=0.1890
+ $X2=0.1620 $Y2=0.1890
r53 30 47 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1890 $X2=0.1890 $Y2=0.1665
r54 30 50 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1890 $X2=0.1755 $Y2=0.1890
r55 24 31 1.49895 $w=1.95333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1485 $X2=0.1890 $Y2=0.1350
r56 24 47 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1485 $X2=0.1890 $Y2=0.1665
r57 31 46 2.6649 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1705 $Y2=0.1350
r58 45 46 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.1545
+ $Y=0.1350 $X2=0.1705 $Y2=0.1350
r59 44 45 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1455
+ $Y=0.1350 $X2=0.1545 $Y2=0.1350
r60 23 44 1.16595 $w=1.3e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1405
+ $Y=0.1350 $X2=0.1455 $Y2=0.1350
r61 42 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1555 $Y=0.1350
+ $X2=0.1545 $Y2=0.1350
r62 41 42 4.72579 $w=1.53e-08 $l=8e-09 $layer=LIG $thickness=4.8e-08 $X=0.1475
+ $Y=0.1350 $X2=0.1555 $Y2=0.1350
r63 39 41 1.73797 $w=1.72143e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1440 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r64 1 39 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.1340
+ $Y=0.1350 $X2=0.1440 $Y2=0.1350
r65 14 1 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1340 $Y2=0.1350
r66 14 41 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r67 7 18 1e-05
r68 6 17 1e-05
.ends

.subckt PM_DHLx3_ASAP7_75t_R%CLKB VSS 9 45 47 13 4 3 12 10 18 11 15 14 1 17 16
c1 1 VSS 9.50386e-20
c2 3 VSS 0.00708318f
c3 4 VSS 0.00720007f
c4 9 VSS 0.00452865f
c5 10 VSS 0.00608167f
c6 11 VSS 0.00602585f
c7 12 VSS 0.0097307f
c8 13 VSS 0.0083787f
c9 14 VSS 0.00628336f
c10 15 VSS 0.000696244f
c11 16 VSS 0.00356348f
c12 17 VSS 0.00307916f
c13 18 VSS 0.00518305f
r1 11 4 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1600 $Y2=0.2160
r2 47 11 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r3 10 3 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1600 $Y2=0.0540
r4 45 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r5 4 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r6 3 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r7 42 43 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1845 $Y2=0.2340
r8 13 17 4.75866 $w=1.41702e-08 $l=2.72259e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.2340 $X2=0.2430 $Y2=0.2305
r9 13 43 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.1845 $Y2=0.2340
r10 39 40 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1845 $Y2=0.0360
r11 12 16 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.0360 $X2=0.2430 $Y2=0.0360
r12 12 40 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.1845 $Y2=0.0360
r13 17 36 3.70931 $w=1.44474e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.2305 $X2=0.2430 $Y2=0.2115
r14 16 34 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0360 $X2=0.2430 $Y2=0.0630
r15 35 36 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1890 $X2=0.2430 $Y2=0.2115
r16 33 34 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0990 $X2=0.2430 $Y2=0.0630
r17 32 33 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1215 $X2=0.2430 $Y2=0.0990
r18 31 35 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1710 $X2=0.2430 $Y2=0.1890
r19 30 31 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1530 $X2=0.2430 $Y2=0.1710
r20 14 30 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1530
r21 14 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1215
r22 28 29 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1530 $X2=0.4050 $Y2=0.1530
r23 27 28 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1530 $X2=0.3240 $Y2=0.1530
r24 27 30 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.2430 $Y=0.1530
+ $X2=0.2430 $Y2=0.1530
r25 18 27 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.2315
+ $Y=0.1530 $X2=0.2430 $Y2=0.1530
r26 25 29 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4050 $Y=0.1530
+ $X2=0.4050 $Y2=0.1530
r27 24 25 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1435 $X2=0.4050 $Y2=0.1530
r28 23 24 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1340 $X2=0.4050 $Y2=0.1435
r29 15 23 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1155 $X2=0.4050 $Y2=0.1340
r30 9 1 5.63117 $w=1.26721e-07 $l=3e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4050 $Y2=0.1320
r31 1 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1320
+ $X2=0.4050 $Y2=0.1340
.ends


*
.SUBCKT DHLx3_ASAP7_75t_R VSS VDD CLK D Q
*
* VSS VSS
* VDD VDD
* CLK CLK
* D D
* Q Q
*
*

MM0 N_MM0_d N_MM0_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2 N_MM2_d N_MM13_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM10_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM6 N_MM6_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM24 N_MM24_d N_MM25_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@3 N_MM24@3_d N_MM25@3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@2 N_MM24@2_d N_MM25@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM12 N_MM12_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM13 N_MM13_d N_MM13_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM25 N_MM25_d N_MM25_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@3 N_MM25@3_d N_MM25@3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@2 N_MM25@2_d N_MM25@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "DHLx3_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "DHLx3_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_DHLx3_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_DHLx3_ASAP7_75t_R%noxref_18
cc_1 N_noxref_18_1 N_MM3_g 0.00135249f
cc_2 N_noxref_18_1 N_CLKB_10 0.000793088f
cc_3 N_noxref_18_1 N_noxref_16_1 0.00768304f
cc_4 N_noxref_18_1 N_noxref_17_1 0.000465156f
x_PM_DHLx3_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_DHLx3_ASAP7_75t_R%noxref_19
cc_5 N_noxref_19_1 N_MM3_g 0.00136187f
cc_6 N_noxref_19_1 N_CLKB_11 0.000740554f
cc_7 N_noxref_19_1 N_noxref_16_1 0.000464293f
cc_8 N_noxref_19_1 N_noxref_17_1 0.00771233f
cc_9 N_noxref_19_1 N_noxref_18_1 0.00123472f
x_PM_DHLx3_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_DHLx3_ASAP7_75t_R%noxref_15
cc_10 N_noxref_15_1 N_MM0_g 0.00366985f
cc_11 N_noxref_15_1 N_CLKN_29 5.51166e-20
cc_12 N_noxref_15_1 N_CLKN_20 8.02379e-20
cc_13 N_noxref_15_1 N_CLKN_28 9.05015e-20
cc_14 N_noxref_15_1 N_CLKN_19 0.000271079f
cc_15 N_noxref_15_1 N_CLKN_7 0.000434691f
cc_16 N_noxref_15_1 N_CLKN_18 0.0276118f
cc_17 N_noxref_15_1 N_noxref_14_1 0.00203831f
x_PM_DHLx3_ASAP7_75t_R%PD3 VSS N_MM9_s N_MM8_d N_PD3_1 PM_DHLx3_ASAP7_75t_R%PD3
cc_18 N_PD3_1 N_MM9_g 0.00776298f
cc_19 N_PD3_1 N_MM11_g 0.00777159f
x_PM_DHLx3_ASAP7_75t_R%CLK VSS CLK N_MM0_g N_CLK_8 N_CLK_6 N_CLK_1 N_CLK_4
+ N_CLK_7 N_CLK_5 PM_DHLx3_ASAP7_75t_R%CLK
x_PM_DHLx3_ASAP7_75t_R%PU1 VSS N_MM3_d N_MM1_s N_PU1_1 PM_DHLx3_ASAP7_75t_R%PU1
cc_20 N_PU1_1 N_MM1_g 0.0170374f
cc_21 N_PU1_1 N_MM3_g 0.017165f
x_PM_DHLx3_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_DHLx3_ASAP7_75t_R%noxref_14
cc_22 N_noxref_14_1 N_MM0_g 0.00370419f
cc_23 N_noxref_14_1 N_CLKN_7 4.28898e-20
cc_24 N_noxref_14_1 N_CLKN_27 5.94188e-20
cc_25 N_noxref_14_1 N_CLKN_19 0.000381583f
cc_26 N_noxref_14_1 N_CLKN_6 0.000504536f
cc_27 N_noxref_14_1 N_CLKN_17 0.0276106f
x_PM_DHLx3_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_DHLx3_ASAP7_75t_R%noxref_16
cc_28 N_noxref_16_1 N_CLKN_1 0.000393237f
cc_29 N_noxref_16_1 N_MM13_g 0.00358831f
cc_30 N_noxref_16_1 N_CLKB_10 0.0274044f
x_PM_DHLx3_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_DHLx3_ASAP7_75t_R%noxref_17
cc_31 N_noxref_17_1 N_CLKN_1 0.000392917f
cc_32 N_noxref_17_1 N_MM13_g 0.0036618f
cc_33 N_noxref_17_1 N_CLKB_11 0.027371f
cc_34 N_noxref_17_1 N_noxref_16_1 0.001432f
x_PM_DHLx3_ASAP7_75t_R%D VSS D N_MM3_g N_D_4 N_D_1 N_D_5 PM_DHLx3_ASAP7_75t_R%D
cc_35 N_D_4 N_CLKN_32 0.000452369f
cc_36 N_D_4 N_CLKN_33 0.000837762f
cc_37 N_D_1 N_CLKN_2 0.00220084f
cc_38 N_MM3_g N_MM1_g 0.00503351f
cc_39 N_D_4 N_CLKN_25 0.00556126f
x_PM_DHLx3_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_DHLx3_ASAP7_75t_R%noxref_21
cc_40 N_noxref_21_1 N_CLKN_8 0.00287403f
cc_41 N_noxref_21_1 N_NET29_11 0.0163163f
cc_42 N_noxref_21_1 N_MM7_g 0.00527724f
cc_43 N_noxref_21_1 N_Q_15 0.000572503f
cc_44 N_noxref_21_1 N_noxref_20_1 0.00148364f
x_PM_DHLx3_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_DHLx3_ASAP7_75t_R%noxref_20
cc_45 N_noxref_20_1 N_NET29_10 0.016998f
cc_46 N_noxref_20_1 N_MH_1 0.000178501f
cc_47 N_noxref_20_1 N_MM7_g 0.00567552f
cc_48 N_noxref_20_1 N_Q_13 0.000751728f
x_PM_DHLx3_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_DHLx3_ASAP7_75t_R%noxref_23
cc_49 N_noxref_23_1 N_CLKN_8 0.000593167f
cc_50 N_noxref_23_1 N_MM25_g 0.00155923f
cc_51 N_noxref_23_1 N_Q_15 0.0366547f
cc_52 N_noxref_23_1 N_noxref_20_1 0.000462944f
cc_53 N_noxref_23_1 N_noxref_21_1 0.00759023f
cc_54 N_noxref_23_1 N_noxref_22_1 0.00122988f
x_PM_DHLx3_ASAP7_75t_R%NET29 VSS N_MM11_g N_MM6_d N_MM7_d N_NET29_4 N_NET29_11
+ N_NET29_16 N_NET29_1 N_NET29_14 N_NET29_3 N_NET29_13 N_NET29_15 N_NET29_10
+ N_NET29_12 N_NET29_17 PM_DHLx3_ASAP7_75t_R%NET29
cc_55 N_MM11_g N_CLKN_3 0.000144457f
cc_56 N_MM11_g N_CLKN_8 0.00481684f
cc_57 N_MM11_g N_CLKN_33 0.000214372f
cc_58 N_MM11_g N_CLKN_26 0.000296527f
cc_59 N_NET29_4 N_CLKN_8 0.00118961f
cc_60 N_NET29_11 N_CLKN_8 0.000382932f
cc_61 N_NET29_16 N_CLKN_8 0.000414079f
cc_62 N_NET29_1 N_MM9_g 0.000424681f
cc_63 N_NET29_14 N_CLKN_8 0.00132055f
cc_64 N_MM11_g N_MM9_g 0.0144087f
x_PM_DHLx3_ASAP7_75t_R%PD2 VSS N_MM10_s N_MM11_d N_PD2_4 N_PD2_5 N_PD2_1
+ PM_DHLx3_ASAP7_75t_R%PD2
cc_65 N_PD2_4 N_CLKN_8 0.000144545f
cc_66 N_PD2_5 N_CLKN_8 0.00111091f
cc_67 N_PD2_1 N_CLKN_3 0.00118169f
cc_68 N_PD2_1 N_MM9_g 0.00232189f
cc_69 N_PD2_5 N_MM9_g 0.0073728f
cc_70 N_PD2_4 N_MM9_g 0.0238641f
cc_71 N_PD2_4 N_MM10_g 0.0149164f
cc_72 N_PD2_5 N_MM11_g 0.0147669f
cc_73 N_PD2_1 N_MH_21 0.000617187f
cc_74 N_PD2_1 N_MH_23 0.000419733f
cc_75 N_PD2_1 N_MH_26 0.000419858f
cc_76 N_PD2_4 N_MH_9 0.000608737f
cc_77 N_PD2_1 N_MH_33 0.00211627f
x_PM_DHLx3_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_DHLx3_ASAP7_75t_R%noxref_24
cc_78 N_noxref_24_1 N_MM25@2_g 0.00151506f
cc_79 N_noxref_24_1 N_Q_14 0.000804127f
x_PM_DHLx3_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_DHLx3_ASAP7_75t_R%noxref_25
cc_80 N_noxref_25_1 N_MM25@2_g 0.00151544f
cc_81 N_noxref_25_1 N_Q_16 0.000815229f
cc_82 N_noxref_25_1 N_noxref_24_1 0.00175251f
x_PM_DHLx3_ASAP7_75t_R%PD1 VSS N_MM5_d N_MM4_s N_PD1_4 N_PD1_5 N_PD1_1
+ PM_DHLx3_ASAP7_75t_R%PD1
cc_83 N_PD1_4 N_CLKN_25 0.000466814f
cc_84 N_PD1_4 N_CLKN_2 0.00239552f
cc_85 N_PD1_4 N_MM1_g 0.0737897f
cc_86 N_PD1_4 N_D_1 0.000646625f
cc_87 N_PD1_4 N_D_4 0.0007279f
cc_88 N_PD1_4 N_MM3_g 0.0358929f
cc_89 N_PD1_5 N_CLKB_1 0.000656526f
cc_90 N_PD1_5 N_MM10_g 0.0348353f
cc_91 N_PD1_1 N_MH_25 9.28656e-20
cc_92 N_PD1_1 N_MH_24 0.000158605f
cc_93 N_PD1_1 N_MH_10 0.00139023f
cc_94 N_PD1_1 N_MH_19 0.00311508f
x_PM_DHLx3_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_DHLx3_ASAP7_75t_R%noxref_22
cc_95 N_noxref_22_1 N_NET29_10 0.000560806f
cc_96 N_noxref_22_1 N_MM25_g 0.00163602f
cc_97 N_noxref_22_1 N_Q_13 0.0364275f
cc_98 N_noxref_22_1 N_noxref_20_1 0.00775603f
cc_99 N_noxref_22_1 N_noxref_21_1 0.000454652f
x_PM_DHLx3_ASAP7_75t_R%Q VSS Q N_MM24_d N_MM24@3_d N_MM24@2_d N_MM25@3_d
+ N_MM25@2_d N_MM25_d N_Q_1 N_Q_18 N_Q_17 N_Q_2 N_Q_14 N_Q_3 N_Q_15 N_Q_13
+ N_Q_19 N_Q_4 N_Q_16 PM_DHLx3_ASAP7_75t_R%Q
cc_100 N_Q_1 N_NET29_14 0.000446362f
cc_101 N_Q_18 N_NET29_16 0.000515456f
cc_102 N_Q_17 N_NET29_17 0.000571548f
cc_103 N_Q_2 N_NET29_14 0.00241576f
cc_104 N_Q_14 N_MM25_g 0.00010294f
cc_105 N_Q_14 N_MH_30 0.000110774f
cc_106 N_Q_14 N_MH_28 0.00013603f
cc_107 N_Q_3 N_MH_29 0.00204449f
cc_108 N_Q_18 N_MH_28 0.000213071f
cc_109 N_Q_18 N_MH_29 0.00240973f
cc_110 N_Q_15 N_MM25_g 0.0156251f
cc_111 N_Q_13 N_MM25_g 0.0525119f
cc_112 N_Q_19 N_MH_30 0.00628853f
cc_113 N_Q_4 N_MH_3 0.000520345f
cc_114 N_Q_2 N_MH_2 0.000693799f
cc_115 N_Q_4 N_MH_4 0.000775026f
cc_116 N_Q_16 N_MM25@3_g 0.0307599f
cc_117 N_Q_16 N_MH_4 0.00130616f
cc_118 N_Q_2 N_MM25_g 0.00133618f
cc_119 N_Q_16 N_MH_3 0.00141158f
cc_120 N_Q_1 N_MM25_g 0.00143842f
cc_121 N_Q_15 N_MH_2 0.00175405f
cc_122 N_Q_1 N_MH_28 0.0019836f
cc_123 N_Q_18 N_MH_34 0.00209927f
cc_124 N_Q_4 N_MM25@3_g 0.00213157f
cc_125 N_Q_3 N_MM25@3_g 0.00218407f
cc_126 N_Q_17 N_MH_29 0.00234002f
cc_127 N_Q_14 N_MM25@2_g 0.0370214f
cc_128 N_Q_14 N_MM25@3_g 0.068116f
x_PM_DHLx3_ASAP7_75t_R%MH VSS N_MM7_g N_MM25_g N_MM25@3_g N_MM25@2_g N_MM4_d
+ N_MM9_d N_MM1_d N_MM10_d N_MH_23 N_MH_32 N_MH_22 N_MH_20 N_MH_9 N_MH_25
+ N_MH_21 N_MH_33 N_MH_1 N_MH_26 N_MH_10 N_MH_34 N_MH_27 N_MH_19 N_MH_24
+ N_MH_28 N_MH_2 N_MH_31 N_MH_30 N_MH_29 N_MH_3 N_MH_4 PM_DHLx3_ASAP7_75t_R%MH
cc_129 N_MH_23 N_CLKN_25 0.000127792f
cc_130 N_MH_32 N_CLKN_26 0.00013598f
cc_131 N_MH_22 N_MM1_g 0.000159182f
cc_132 N_MH_20 N_MM9_g 0.000162247f
cc_133 N_MH_9 N_CLKN_2 0.000253141f
cc_134 N_MH_25 N_CLKN_26 0.000256976f
cc_135 N_MH_21 N_MM1_g 0.0346187f
cc_136 N_MH_33 N_CLKN_26 0.000334588f
cc_137 N_MH_9 N_CLKN_32 0.000354108f
cc_138 N_MH_9 N_CLKN_25 0.000521854f
cc_139 N_MH_1 N_CLKN_8 0.00176768f
cc_140 N_MH_26 N_CLKN_33 0.000589348f
cc_141 N_MH_10 N_MM9_g 0.000645104f
cc_142 N_MH_34 N_CLKN_26 0.000647698f
cc_143 N_MH_27 N_CLKN_8 0.00065136f
cc_144 N_MH_21 N_CLKN_2 0.00073975f
cc_145 N_MH_26 N_CLKN_3 0.000916226f
cc_146 N_MH_9 N_MM1_g 0.0019236f
cc_147 N_MH_27 N_CLKN_26 0.00205625f
cc_148 N_MH_23 N_CLKN_32 0.00369075f
cc_149 N_MH_26 N_CLKN_26 0.0046539f
cc_150 N_MH_34 N_CLKN_8 0.0047451f
cc_151 N_MH_23 N_CLKN_33 0.00589859f
cc_152 N_MM7_g N_CLKN_8 0.00627307f
cc_153 N_MH_19 N_MM9_g 0.036934f
cc_154 N_MH_27 N_MM10_g 9.53223e-20
cc_155 N_MH_20 N_MM10_g 0.000145946f
cc_156 N_MH_22 N_MM10_g 0.000164091f
cc_157 N_MH_24 N_CLKB_15 0.000234368f
cc_158 N_MH_23 N_CLKB_15 0.000283778f
cc_159 N_MH_21 N_MM10_g 0.0167289f
cc_160 N_MH_34 N_CLKB_18 0.000760223f
cc_161 N_MH_10 N_CLKB_1 0.000788114f
cc_162 N_MH_25 N_CLKB_15 0.000795124f
cc_163 N_MH_26 N_CLKB_15 0.00173476f
cc_164 N_MH_23 N_CLKB_18 0.000933637f
cc_165 N_MH_10 N_MM10_g 0.00113235f
cc_166 N_MH_9 N_MM10_g 0.00116044f
cc_167 N_MH_19 N_CLKB_1 0.00168729f
cc_168 N_MH_32 N_CLKB_15 0.00305788f
cc_169 N_MH_19 N_MM10_g 0.0534443f
cc_170 N_MH_32 N_MM11_g 6.00202e-20
cc_171 N_MH_24 N_MM11_g 6.09855e-20
cc_172 N_MH_28 N_MM11_g 7.37879e-20
cc_173 N_MH_2 N_MM11_g 9.98996e-20
cc_174 N_MH_19 N_MM11_g 0.000162457f
cc_175 N_MH_27 N_MM11_g 0.000163183f
cc_176 N_MM7_g N_NET29_11 0.00669391f
cc_177 N_MM7_g N_NET29_3 0.000355529f
cc_178 N_MH_34 N_NET29_16 0.000410672f
cc_179 N_MH_10 N_NET29_1 0.000453379f
cc_180 N_MH_28 N_NET29_14 0.000458242f
cc_181 N_MH_27 N_NET29_13 0.00068194f
cc_182 N_MH_1 N_NET29_14 0.000801356f
cc_183 N_MH_27 N_NET29_1 0.000919156f
cc_184 N_MH_1 N_MM11_g 0.000931781f
cc_185 N_MH_31 N_NET29_15 0.000972126f
cc_186 N_MM7_g N_NET29_1 0.00108469f
cc_187 N_MM7_g N_NET29_10 0.00650297f
cc_188 N_MH_34 N_NET29_14 0.00262358f
cc_189 N_MH_27 N_NET29_12 0.00303111f
cc_190 N_MH_25 N_NET29_12 0.00356398f
cc_191 N_MH_27 N_NET29_14 0.00404456f
cc_192 N_MM7_g N_MM11_g 0.0290876f
x_PM_DHLx3_ASAP7_75t_R%CLKN VSS N_MM13_g N_MM1_g N_MM9_g N_MM0_d N_MM12_d
+ N_CLKN_24 N_CLKN_31 N_CLKN_28 N_CLKN_30 N_CLKN_7 N_CLKN_6 N_CLKN_18 N_CLKN_17
+ N_CLKN_1 N_CLKN_22 N_CLKN_19 N_CLKN_23 N_CLKN_33 N_CLKN_21 N_CLKN_32 N_CLKN_2
+ N_CLKN_25 N_CLKN_8 N_CLKN_3 N_CLKN_26 N_CLKN_27 N_CLKN_29 N_CLKN_20
+ PM_DHLx3_ASAP7_75t_R%CLKN
cc_193 N_CLKN_24 N_MM0_g 8.56612e-20
cc_194 N_CLKN_31 N_MM0_g 0.00012494f
cc_195 N_CLKN_28 N_MM0_g 0.000185001f
cc_196 N_CLKN_30 N_MM0_g 0.000187207f
cc_197 N_CLKN_7 N_MM0_g 0.00105024f
cc_198 N_CLKN_6 N_MM0_g 0.00114354f
cc_199 N_CLKN_18 N_MM0_g 0.0112134f
cc_200 N_CLKN_17 N_MM0_g 0.0112205f
cc_201 N_CLKN_1 N_CLK_8 0.000430464f
cc_202 N_CLKN_22 N_CLK_6 0.000666503f
cc_203 N_CLKN_1 N_CLK_1 0.00340882f
cc_204 N_CLKN_19 N_CLK_4 0.000993062f
cc_205 N_CLKN_23 N_CLK_8 0.00127749f
cc_206 N_CLKN_23 N_CLK_7 0.00139399f
cc_207 N_CLKN_30 N_CLK_8 0.00151226f
cc_208 N_CLKN_33 N_CLK_6 0.00176626f
cc_209 N_CLKN_21 N_CLK_5 0.00185753f
cc_210 N_CLKN_30 N_CLK_6 0.00233153f
cc_211 N_CLKN_28 N_CLK_8 0.00287257f
cc_212 N_CLKN_19 N_CLK_7 0.00297601f
cc_213 N_MM13_g N_MM0_g 0.0350987f
x_PM_DHLx3_ASAP7_75t_R%CLKB VSS N_MM10_g N_MM2_d N_MM13_d N_CLKB_13 N_CLKB_4
+ N_CLKB_3 N_CLKB_12 N_CLKB_10 N_CLKB_18 N_CLKB_11 N_CLKB_15 N_CLKB_14 N_CLKB_1
+ N_CLKB_17 N_CLKB_16 PM_DHLx3_ASAP7_75t_R%CLKB
cc_214 N_CLKB_13 N_CLK_5 0.000181951f
cc_215 N_CLKB_4 N_CLK_5 0.000198639f
cc_216 N_CLKB_3 N_CLK_5 0.000266327f
cc_217 N_CLKB_13 N_CLK_6 0.00105956f
cc_218 N_CLKB_12 N_CLK_5 0.00269212f
cc_219 N_CLKB_10 N_CLKN_19 5.85679e-20
cc_220 N_CLKB_10 N_CLKN_8 0.000112543f
cc_221 N_CLKB_10 N_CLKN_30 0.000240245f
cc_222 N_CLKB_4 N_CLKN_30 0.000286722f
cc_223 N_CLKB_13 N_CLKN_30 0.00513698f
cc_224 N_CLKB_18 N_CLKN_25 0.000389596f
cc_225 N_CLKB_11 N_MM13_g 0.0112874f
cc_226 N_CLKB_4 N_CLKN_1 0.000405695f
cc_227 N_CLKB_12 N_CLKN_31 0.000473999f
cc_228 N_CLKB_15 N_CLKN_32 0.000486429f
cc_229 N_CLKB_14 N_CLKN_23 0.000587202f
cc_230 N_MM10_g N_CLKN_3 0.000615758f
cc_231 N_CLKB_15 N_CLKN_33 0.000680446f
cc_232 N_CLKB_3 N_MM13_g 0.000761329f
cc_233 N_CLKB_1 N_CLKN_2 0.00220715f
cc_234 N_CLKB_11 N_CLKN_1 0.000935649f
cc_235 N_CLKB_14 N_CLKN_33 0.000943698f
cc_236 N_CLKB_14 N_CLKN_24 0.00109687f
cc_237 N_CLKB_4 N_MM13_g 0.0011332f
cc_238 N_CLKB_15 N_CLKN_25 0.00365005f
cc_239 N_MM10_g N_MM9_g 0.00368403f
cc_240 N_CLKB_14 N_CLKN_31 0.00402222f
cc_241 N_MM10_g N_MM1_g 0.00705092f
cc_242 N_CLKB_18 N_CLKN_33 0.0194752f
cc_243 N_CLKB_10 N_MM13_g 0.0389974f
cc_244 N_CLKB_17 N_D_4 0.000365506f
cc_245 N_CLKB_18 N_D_4 0.00104672f
cc_246 N_CLKB_16 N_D_5 0.00108937f
cc_247 N_CLKB_14 N_D_4 0.00861212f
*END of DHLx3_ASAP7_75t_R.pxi
.ENDS
** Design:	DLLx1_ASAP7_75t_R
* Created:	"Fri Aug 17 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "DLLx1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "DLLx1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_DLLx1_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.0041966f
.ends

.subckt PM_DLLx1_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00416324f
.ends

.subckt PM_DLLx1_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.00453477f
.ends

.subckt PM_DLLx1_ASAP7_75t_R%Q VSS 19 14 27 7 2 11 1 8 10
c1 1 VSS 0.00802336f
c2 2 VSS 0.00852081f
c3 7 VSS 0.00375458f
c4 8 VSS 0.00374769f
c5 9 VSS 0.00464961f
c6 10 VSS 0.00362886f
c7 11 VSS 0.00568515f
c8 12 VSS 0.00310349f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7415 $Y=0.2025 $X2=0.7540 $Y2=0.2025
r2 27 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.2025 $X2=0.7415 $Y2=0.2025
r3 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7560 $Y=0.2025
+ $X2=0.7560 $Y2=0.2340
r4 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.2340 $X2=0.7695 $Y2=0.2340
r5 11 22 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7830 $Y=0.2340 $X2=0.7830 $Y2=0.2125
r6 11 25 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7830 $Y=0.2340 $X2=0.7695 $Y2=0.2340
r7 21 22 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1530 $X2=0.7830 $Y2=0.2125
r8 20 21 13.8165 $w=1.3e-08 $l=5.93e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.0937 $X2=0.7830 $Y2=0.1530
r9 19 20 2.97317 $w=1.3e-08 $l=1.27e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.0810 $X2=0.7830 $Y2=0.0937
r10 19 10 4.25571 $w=1.3e-08 $l=1.83e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.0810 $X2=0.7830 $Y2=0.0627
r11 10 12 4.58871 $w=1.62972e-08 $l=2.67e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7830 $Y=0.0627 $X2=0.7830 $Y2=0.0360
r12 12 18 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7830 $Y=0.0360 $X2=0.7695 $Y2=0.0360
r13 17 18 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.0360 $X2=0.7695 $Y2=0.0360
r14 16 17 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.7445
+ $Y=0.0360 $X2=0.7560 $Y2=0.0360
r15 9 16 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.7400
+ $Y=0.0360 $X2=0.7445 $Y2=0.0360
r16 1 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7560 $Y=0.0675
+ $X2=0.7560 $Y2=0.0360
r17 7 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7415 $Y=0.0675 $X2=0.7540 $Y2=0.0675
r18 14 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.0675 $X2=0.7415 $Y2=0.0675
.ends

.subckt PM_DLLx1_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.0417514f
.ends

.subckt PM_DLLx1_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.00478329f
.ends

.subckt PM_DLLx1_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.00462738f
.ends

.subckt PM_DLLx1_ASAP7_75t_R%PD3 VSS 2 4 1
c1 1 VSS 0.000930846f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0405 $X2=0.4905 $Y2=0.0405
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0405 $X2=0.4735 $Y2=0.0405
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4735 $Y=0.0405 $X2=0.4905 $Y2=0.0405
.ends

.subckt PM_DLLx1_ASAP7_75t_R%PU1 VSS 2 4 1
c1 1 VSS 0.000968213f
r1 4 3 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3365 $Y2=0.2025
r2 2 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3195 $Y2=0.2025
r3 1 3 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3195 $Y=0.2025 $X2=0.3365 $Y2=0.2025
.ends

.subckt PM_DLLx1_ASAP7_75t_R%PD1 VSS 7 10 5 4 1
c1 1 VSS 0.00934602f
c2 4 VSS 0.00316954f
c3 5 VSS 0.00186607f
r1 10 9 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r2 8 9 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r3 5 8 0.123457 $w=8.1e-08 $l=1e-08 $layer=N_src_drn $thickness=1e-09 $X=0.3780
+ $Y=0.0675 $X2=0.3880 $Y2=0.0675
r4 4 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3220 $Y2=0.0675
r5 7 4 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r6 1 5 1e-05
.ends

.subckt PM_DLLx1_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.0417915f
.ends

.subckt PM_DLLx1_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.0418419f
.ends

.subckt PM_DLLx1_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.00469065f
.ends

.subckt PM_DLLx1_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.0046708f
.ends

.subckt PM_DLLx1_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.00365655f
.ends

.subckt PM_DLLx1_ASAP7_75t_R%PD2 VSS 7 13 4 5 1
c1 1 VSS 0.00713671f
c2 4 VSS 0.00187869f
c3 5 VSS 0.00234016f
r1 13 12 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r2 5 12 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4880 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r3 10 5 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4725
+ $Y=0.2295 $X2=0.4860 $Y2=0.2295
r4 9 10 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4590
+ $Y=0.2295 $X2=0.4725 $Y2=0.2295
r5 8 9 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4455
+ $Y=0.2295 $X2=0.4590 $Y2=0.2295
r6 1 8 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4320
+ $Y=0.2295 $X2=0.4455 $Y2=0.2295
r7 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2295 $X2=0.4300 $Y2=0.2295
r8 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2295 $X2=0.4175 $Y2=0.2295
.ends

.subckt PM_DLLx1_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.041942f
.ends

.subckt PM_DLLx1_ASAP7_75t_R%MH VSS 11 12 63 67 71 75 21 5 16 18 15 24 26 19 20
+ 17 6 13 14 25 1 2 22 23
c1 1 VSS 0.000457238f
c2 2 VSS 0.00405262f
c3 5 VSS 0.00619103f
c4 6 VSS 0.00503663f
c5 11 VSS 0.0369431f
c6 12 VSS 0.0802329f
c7 13 VSS 0.00308436f
c8 14 VSS 0.000453722f
c9 15 VSS 0.00355021f
c10 16 VSS 0.00043915f
c11 17 VSS 0.00773417f
c12 18 VSS 0.00374353f
c13 19 VSS 0.00107515f
c14 20 VSS 0.000688671f
c15 21 VSS 0.00052891f
c16 22 VSS 0.00382404f
c17 23 VSS 0.00247179f
c18 24 VSS 2.61715e-20
c19 25 VSS 0.00243948f
c20 26 VSS 0.00709019f
r1 75 74 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r2 73 74 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r3 15 73 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3760 $Y=0.2295 $X2=0.3880 $Y2=0.2295
r4 16 15 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2295 $X2=0.3760 $Y2=0.2295
r5 69 70 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r6 71 69 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.1890 $X2=0.3635 $Y2=0.1890
r7 15 70 0.185185 $w=5.4e-08 $l=1e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r8 67 66 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r9 65 66 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4420 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r10 6 65 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4300 $Y=0.0405 $X2=0.4420 $Y2=0.0405
r11 14 6 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0405 $X2=0.4300 $Y2=0.0405
r12 13 6 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0810 $X2=0.4300 $Y2=0.0810
r13 63 13 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0810 $X2=0.4175 $Y2=0.0810
r14 59 15 15.0298 $w=2.02e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.3780 $Y=0.2045 $X2=0.3780 $Y2=0.1790
r15 5 52 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2295
+ $X2=0.3780 $Y2=0.2340
r16 5 59 14.7351 $w=2.02e-08 $l=2.5e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.3780 $Y=0.2295 $X2=0.3780 $Y2=0.2045
r17 2 48 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7290 $Y=0.1360
+ $X2=0.7290 $Y2=0.1445
r18 12 2 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=0.7290
+ $Y=0.1350 $X2=0.7290 $Y2=0.1360
r19 6 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0405
+ $X2=0.4320 $Y2=0.0360
r20 52 53 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r21 50 53 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r22 17 25 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4320 $Y=0.2340 $X2=0.4590 $Y2=0.2340
r23 17 50 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4050 $Y2=0.2340
r24 22 48 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1165 $X2=0.7290 $Y2=0.1445
r25 18 23 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4320 $Y=0.0360 $X2=0.4590 $Y2=0.0360
r26 25 43 3.01468 $w=1.741e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4590 $Y2=0.2140
r27 46 48 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.7290 $Y=0.1530
+ $X2=0.7290 $Y2=0.1445
r28 45 46 24.6015 $w=1.3e-08 $l=1.055e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.6235 $Y=0.1530 $X2=0.7290 $Y2=0.1530
r29 44 45 29.3819 $w=1.3e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.4975
+ $Y=0.1530 $X2=0.6235 $Y2=0.1530
r30 26 44 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M2 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1530 $X2=0.4975 $Y2=0.1530
r31 26 39 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4590 $Y=0.1530
+ $X2=0.4590 $Y2=0.1530
r32 23 38 6.51253 $w=1.552e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4590 $Y2=0.0710
r33 42 43 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2015 $X2=0.4590 $Y2=0.2140
r34 41 42 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1825 $X2=0.4590 $Y2=0.2015
r35 40 41 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1635 $X2=0.4590 $Y2=0.1825
r36 39 40 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1530 $X2=0.4590 $Y2=0.1635
r37 20 39 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1420 $X2=0.4590 $Y2=0.1530
r38 20 24 1.38478 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1420 $X2=0.4590 $Y2=0.1310
r39 37 38 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1015 $X2=0.4590 $Y2=0.0710
r40 19 24 2.78392 $w=1.56471e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1140 $X2=0.4590 $Y2=0.1310
r41 19 37 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1140 $X2=0.4590 $Y2=0.1015
r42 24 36 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1310 $X2=0.4860 $Y2=0.1310
r43 35 36 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1310 $X2=0.4860 $Y2=0.1310
r44 21 33 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.5395
+ $Y=0.1310 $X2=0.5660 $Y2=0.1310
r45 21 35 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.5395
+ $Y=0.1310 $X2=0.5130 $Y2=0.1310
r46 1 30 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.5670
+ $Y=0.1310 $X2=0.5670 $Y2=0.1310
r47 1 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1310
+ $X2=0.5660 $Y2=0.1310
r48 11 30 0.314665 $w=2.27e-07 $l=4e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5670 $Y=0.1350 $X2=0.5670 $Y2=0.1310
.ends

.subckt PM_DLLx1_ASAP7_75t_R%CLK VSS 11 3 8 6 1 7 5 4
c1 1 VSS 0.00254732f
c2 3 VSS 0.0597268f
c3 4 VSS 0.000795114f
c4 5 VSS 0.0042528f
c5 6 VSS 0.00412861f
c6 7 VSS 0.00190601f
c7 8 VSS 0.00179212f
r1 6 17 2.40741 $w=2.45e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.1980 $X2=0.1080 $Y2=0.1710
r2 5 15 4.50612 $w=2.06667e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0630 $X2=0.1080 $Y2=0.0990
r3 16 17 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.1710 $X2=0.1080 $Y2=0.1710
r4 8 13 1.35805 $w=2.83333e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1710 $X2=0.0810 $Y2=0.1485
r5 8 16 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1710 $X2=0.0945 $Y2=0.1710
r6 14 15 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.0990 $X2=0.1080 $Y2=0.0990
r7 7 10 0.483592 $w=3.42308e-08 $l=1.87e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0990 $X2=0.0810 $Y2=0.1177
r8 7 14 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0990 $X2=0.0945 $Y2=0.0990
r9 11 12 0.874462 $w=1.3e-08 $l=3.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1227
r10 11 10 0.291487 $w=1.3e-08 $l=1.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1177
r11 4 12 2.85657 $w=1.3e-08 $l=1.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1227
r12 4 13 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1485
r13 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r14 1 4 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_DLLx1_ASAP7_75t_R%D VSS 9 3 4 5 6 1
c1 1 VSS 0.00653833f
c2 3 VSS 0.0833577f
c3 4 VSS 0.00563718f
c4 5 VSS 0.00673646f
c5 6 VSS 0.00728371f
r1 6 13 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.2340 $X2=0.2970 $Y2=0.2140
r2 12 13 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1735 $X2=0.2970 $Y2=0.2140
r3 11 12 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1735
r4 10 11 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1215 $X2=0.2970 $Y2=0.1350
r5 9 10 1.16595 $w=1.3e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1165 $X2=0.2970 $Y2=0.1215
r6 9 8 1.28254 $w=1.3e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1165 $X2=0.2970 $Y2=0.1110
r7 4 8 8.27824 $w=1.3e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0755 $X2=0.2970 $Y2=0.1110
r8 4 5 8.03069 $w=1.41392e-08 $l=3.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0755 $X2=0.2970 $Y2=0.0360
r9 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r10 1 11 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_DLLx1_ASAP7_75t_R%NET085 VSS 9 35 40 16 11 1 4 14 3 13 15 10 12
c1 1 VSS 0.00286952f
c2 3 VSS 0.00597229f
c3 4 VSS 0.00640634f
c4 9 VSS 0.0375167f
c5 10 VSS 0.00332185f
c6 11 VSS 0.00350397f
c7 12 VSS 0.0012605f
c8 13 VSS 0.00828349f
c9 14 VSS 0.00524123f
c10 15 VSS 0.00281197f
c11 16 VSS 0.00614209f
c12 17 VSS 0.00371046f
r1 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2295 $X2=0.5920 $Y2=0.2295
r2 40 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.2295 $X2=0.5795 $Y2=0.2295
r3 4 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2295
+ $X2=0.5940 $Y2=0.2340
r4 37 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.2340 $X2=0.6075 $Y2=0.2340
r5 16 33 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.2340 $X2=0.6210 $Y2=0.2140
r6 16 38 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.2340 $X2=0.6075 $Y2=0.2340
r7 10 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.0405 $X2=0.5920 $Y2=0.0405
r8 35 10 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0405 $X2=0.5795 $Y2=0.0405
r9 32 33 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.2015 $X2=0.6210 $Y2=0.2140
r10 31 32 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1825 $X2=0.6210 $Y2=0.2015
r11 30 31 6.99569 $w=1.3e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1525 $X2=0.6210 $Y2=0.1825
r12 29 30 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1310 $X2=0.6210 $Y2=0.1525
r13 28 29 3.96423 $w=1.3e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1140 $X2=0.6210 $Y2=0.1310
r14 27 28 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1015 $X2=0.6210 $Y2=0.1140
r15 14 17 6.51253 $w=1.552e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.0710 $X2=0.6210 $Y2=0.0360
r16 14 27 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0710 $X2=0.6210 $Y2=0.1015
r17 3 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0405
+ $X2=0.5940 $Y2=0.0360
r18 17 26 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.0360 $X2=0.6075 $Y2=0.0360
r19 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0360 $X2=0.6075 $Y2=0.0360
r20 24 25 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5825
+ $Y=0.0360 $X2=0.5940 $Y2=0.0360
r21 13 15 7.2121 $w=1.41842e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5510 $Y=0.0360 $X2=0.5130 $Y2=0.0360
r22 13 24 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5510
+ $Y=0.0360 $X2=0.5825 $Y2=0.0360
r23 12 22 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0590 $X2=0.5130 $Y2=0.0820
r24 12 15 3.71425 $w=1.68348e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.0590 $X2=0.5130 $Y2=0.0360
r25 1 19 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.5130
+ $Y=0.0820 $X2=0.5130 $Y2=0.0820
r26 1 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.0820
+ $X2=0.5130 $Y2=0.0820
r27 9 19 0.314665 $w=2.27e-07 $l=5.3e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5130 $Y2=0.0820
.ends

.subckt PM_DLLx1_ASAP7_75t_R%CLKN VSS 11 12 67 69 6 5 23 13 14 1 16 18 19 17 27
+ 25 15 21 20 26 2
c1 1 VSS 0.00166069f
c2 2 VSS 7.19883e-20
c3 5 VSS 0.00755988f
c4 6 VSS 0.00760135f
c5 11 VSS 0.0597516f
c6 12 VSS 0.00453872f
c7 13 VSS 0.00566047f
c8 14 VSS 0.00566718f
c9 15 VSS 0.00494268f
c10 16 VSS 0.00318544f
c11 17 VSS 0.00480534f
c12 18 VSS 0.0046017f
c13 19 VSS 0.000423732f
c14 20 VSS 0.000373191f
c15 21 VSS 0.000769385f
c16 22 VSS 0.00361801f
c17 23 VSS 0.00142637f
c18 24 VSS 0.0034594f
c19 25 VSS 0.000792523f
c20 26 VSS 0.000405455f
c21 27 VSS 0.0139294f
r1 69 68 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r2 14 68 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r3 67 66 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r4 13 66 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r5 11 60 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1340 $Y2=0.1350
r6 6 57 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0550 $Y2=0.2340
r7 5 54 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0550 $Y2=0.0360
r8 60 61 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.1340
+ $Y=0.1350 $X2=0.1440 $Y2=0.1350
r9 1 61 1.73797 $w=1.72143e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1475 $Y=0.1350 $X2=0.1440 $Y2=0.1350
r10 1 63 4.72579 $w=1.53e-08 $l=8e-09 $layer=LIG $thickness=4.8e-08 $X=0.1475
+ $Y=0.1350 $X2=0.1555 $Y2=0.1350
r11 56 57 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.2340 $X2=0.0550 $Y2=0.2340
r12 18 56 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0460 $Y2=0.2340
r13 18 24 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0180 $Y2=0.2340
r14 53 54 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.0360 $X2=0.0550 $Y2=0.0360
r15 17 53 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0460 $Y2=0.0360
r16 17 22 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0180 $Y2=0.0360
r17 19 50 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.1545
+ $Y=0.1350 $X2=0.1705 $Y2=0.1350
r18 19 63 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1545 $Y=0.1350
+ $X2=0.1555 $Y2=0.1350
r19 24 48 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.2340 $X2=0.0180 $Y2=0.2070
r20 22 47 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.0360 $X2=0.0180 $Y2=0.0630
r21 25 45 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1980 $X2=0.1890 $Y2=0.1755
r22 26 50 2.6649 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1705 $Y2=0.1350
r23 16 23 3.9134 $w=1.47857e-08 $l=2.25499e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1755 $X2=0.0165 $Y2=0.1530
r24 16 48 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1755 $X2=0.0180 $Y2=0.2070
r25 46 47 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0990 $X2=0.0180 $Y2=0.0630
r26 15 23 3.9134 $w=1.47857e-08 $l=2.25499e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1305 $X2=0.0165 $Y2=0.1530
r27 15 46 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1305 $X2=0.0180 $Y2=0.0990
r28 44 45 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1575 $X2=0.1890 $Y2=0.1755
r29 20 39 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1890 $Y=0.1485
+ $X2=0.1890 $Y2=0.1530
r30 20 44 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1485 $X2=0.1890 $Y2=0.1575
r31 20 26 1.49895 $w=1.95333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1485 $X2=0.1890 $Y2=0.1350
r32 41 42 1.90199 $w=1.38333e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.0255 $Y=0.1530 $X2=0.0345 $Y2=0.1530
r33 23 41 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0165
+ $Y=0.1530 $X2=0.0255 $Y2=0.1530
r34 39 40 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1530 $X2=0.2135 $Y2=0.1530
r35 38 39 18.1888 $w=1.3e-08 $l=7.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.1110
+ $Y=0.1530 $X2=0.1890 $Y2=0.1530
r36 37 38 18.1888 $w=1.3e-08 $l=7.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.0330
+ $Y=0.1530 $X2=0.1110 $Y2=0.1530
r37 37 42 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.0330 $Y=0.1530
+ $X2=0.0345 $Y2=0.1530
r38 27 35 21.5701 $w=1.3e-08 $l=9.25e-08 $layer=M2 $thickness=3.6e-08 $X=0.3125
+ $Y=0.1530 $X2=0.4050 $Y2=0.1530
r39 27 40 23.0858 $w=1.3e-08 $l=9.9e-08 $layer=M2 $thickness=3.6e-08 $X=0.3125
+ $Y=0.1530 $X2=0.2135 $Y2=0.1530
r40 33 35 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4050 $Y=0.1440
+ $X2=0.4050 $Y2=0.1530
r41 21 33 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1160 $X2=0.4050 $Y2=0.1440
r42 12 2 5.63117 $w=1.26721e-07 $l=2e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4050 $Y2=0.1330
r43 2 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1330
+ $X2=0.4050 $Y2=0.1440
r44 6 14 1e-05
r45 5 13 1e-05
.ends

.subckt PM_DLLx1_ASAP7_75t_R%CLKB VSS 12 13 71 73 14 5 17 4 16 21 6 15 19 18 23
+ 2 1 22 20
c1 1 VSS 0.000280591f
c2 2 VSS 9.02939e-20
c3 4 VSS 0.00690983f
c4 5 VSS 0.0072179f
c5 6 VSS 0.00493872f
c6 12 VSS 0.0052636f
c7 13 VSS 0.00507709f
c8 14 VSS 0.00629352f
c9 15 VSS 0.00624923f
c10 16 VSS 0.00927456f
c11 17 VSS 0.00896048f
c12 18 VSS 0.00613713f
c13 19 VSS 0.00119219f
c14 20 VSS 0.00151669f
c15 21 VSS 0.00315481f
c16 22 VSS 0.0030436f
c17 23 VSS 0.0109902f
r1 15 5 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1600 $Y2=0.2160
r2 73 15 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r3 14 4 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1600 $Y2=0.0540
r4 71 14 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r5 5 66 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r6 4 63 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r7 2 54 5.67512 $w=2.4e-08 $l=5e-09 $layer=LISD $thickness=4.02632e-08
+ $X=0.4590 $Y=0.1790 $X2=0.4640 $Y2=0.1790
r8 13 2 2.88446 $w=1.16273e-07 $l=4.4e-08 $layer=LIG $thickness=5.16364e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4590 $Y2=0.1790
r9 66 67 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1845 $Y2=0.2340
r10 17 22 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.2340 $X2=0.2430 $Y2=0.2340
r11 17 67 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.1845 $Y2=0.2340
r12 63 64 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1845 $Y2=0.0360
r13 16 21 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.0360 $X2=0.2430 $Y2=0.0360
r14 16 64 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.1845 $Y2=0.0360
r15 52 54 11.0623 $w=2.14976e-08 $l=2.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4845 $Y=0.1790 $X2=0.4640 $Y2=0.1790
r16 51 52 8.84105 $w=2.02e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4995 $Y=0.1790 $X2=0.4845 $Y2=0.1790
r17 6 49 6.18874 $w=2.02e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5025 $Y=0.1790 $X2=0.5130 $Y2=0.1790
r18 6 51 1.76821 $w=2.02e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.5025
+ $Y=0.1790 $X2=0.4995 $Y2=0.1790
r19 22 46 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2430 $Y2=0.2160
r20 21 43 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0360 $X2=0.2430 $Y2=0.0630
r21 47 49 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5130 $Y=0.1845
+ $X2=0.5130 $Y2=0.1790
r22 20 47 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1680 $X2=0.5130 $Y2=0.1845
r23 45 46 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2025 $X2=0.2430 $Y2=0.2160
r24 44 45 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1935 $X2=0.2430 $Y2=0.2025
r25 42 43 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0990 $X2=0.2430 $Y2=0.0630
r26 41 42 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1215 $X2=0.2430 $Y2=0.0990
r27 40 44 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1845 $X2=0.2430 $Y2=0.1935
r28 18 40 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1530 $X2=0.2430 $Y2=0.1845
r29 18 41 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1530 $X2=0.2430 $Y2=0.1215
r30 38 47 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.5130 $Y=0.1890
+ $X2=0.5130 $Y2=0.1845
r31 37 38 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.4770
+ $Y=0.1890 $X2=0.5130 $Y2=0.1890
r32 36 37 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M2 $thickness=3.6e-08 $X=0.4320
+ $Y=0.1890 $X2=0.4770 $Y2=0.1890
r33 35 36 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M2 $thickness=3.6e-08 $X=0.3870
+ $Y=0.1890 $X2=0.4320 $Y2=0.1890
r34 34 35 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1890 $X2=0.3870 $Y2=0.1890
r35 33 34 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1890 $X2=0.3510 $Y2=0.1890
r36 32 33 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1890 $X2=0.2970 $Y2=0.1890
r37 32 40 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.2430 $Y=0.1890
+ $X2=0.2430 $Y2=0.1845
r38 23 32 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.2315
+ $Y=0.1890 $X2=0.2430 $Y2=0.1890
r39 29 34 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.3510 $Y=0.1890
+ $X2=0.3510 $Y2=0.1890
r40 28 29 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1620 $X2=0.3510 $Y2=0.1890
r41 27 28 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1620
r42 19 27 4.4306 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1160 $X2=0.3510 $Y2=0.1350
r43 12 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r44 1 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
.ends


*
.SUBCKT DLLx1_ASAP7_75t_R VSS VDD CLK D Q
*
* VSS VSS
* VDD VDD
* CLK CLK
* D D
* Q Q
*
*

MM20 N_MM20_d N_MM20_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM23 N_MM23_d N_MM23_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM10_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM6 N_MM6_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM24 N_MM24_d N_MM25_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM21 N_MM21_d N_MM20_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM22 N_MM22_d N_MM23_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM25 N_MM25_d N_MM25_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "DLLx1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "DLLx1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_DLLx1_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_DLLx1_ASAP7_75t_R%noxref_14
cc_1 N_noxref_14_1 N_MM20_g 0.00367791f
cc_2 N_noxref_14_1 N_CLKN_15 0.000315663f
cc_3 N_noxref_14_1 N_CLKN_5 0.000503546f
cc_4 N_noxref_14_1 N_CLKN_13 0.0278695f
x_PM_DLLx1_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_DLLx1_ASAP7_75t_R%noxref_15
cc_5 N_noxref_15_1 N_MM20_g 0.00366547f
cc_6 N_noxref_15_1 N_CLKN_16 0.000199259f
cc_7 N_noxref_15_1 N_CLKN_6 0.000504268f
cc_8 N_noxref_15_1 N_CLKN_14 0.0281017f
cc_9 N_noxref_15_1 N_noxref_14_1 0.00204313f
x_PM_DLLx1_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_DLLx1_ASAP7_75t_R%noxref_25
cc_10 N_noxref_25_1 N_MM25_g 0.00149703f
cc_11 N_noxref_25_1 N_Q_8 0.0385707f
cc_12 N_noxref_25_1 N_noxref_24_1 0.00177936f
x_PM_DLLx1_ASAP7_75t_R%Q VSS Q N_MM24_d N_MM25_d N_Q_7 N_Q_2 N_Q_11 N_Q_1 N_Q_8
+ N_Q_10 PM_DLLx1_ASAP7_75t_R%Q
cc_13 N_Q_7 N_MH_22 0.00134502f
cc_14 N_Q_2 N_MH_2 0.000843473f
cc_15 N_Q_11 N_MH_26 0.000849145f
cc_16 N_Q_1 N_MM25_g 0.001124f
cc_17 N_Q_2 N_MM25_g 0.00138215f
cc_18 N_Q_8 N_MH_2 0.00160109f
cc_19 N_Q_8 N_MM25_g 0.0154802f
cc_20 N_Q_10 N_MH_22 0.006249f
cc_21 N_Q_7 N_MM25_g 0.0545103f
x_PM_DLLx1_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_DLLx1_ASAP7_75t_R%noxref_22
cc_22 N_noxref_22_1 N_NET085_10 0.00056058f
cc_23 N_noxref_22_1 N_MM25_g 0.00160622f
cc_24 N_noxref_22_1 N_noxref_20_1 0.00774799f
cc_25 N_noxref_22_1 N_noxref_21_1 0.000449197f
x_PM_DLLx1_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_DLLx1_ASAP7_75t_R%noxref_24
cc_26 N_noxref_24_1 N_MM25_g 0.00149486f
cc_27 N_noxref_24_1 N_Q_7 0.0383936f
x_PM_DLLx1_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_DLLx1_ASAP7_75t_R%noxref_20
cc_28 N_noxref_20_1 N_NET085_10 0.0170321f
cc_29 N_noxref_20_1 N_MM7_g 0.00583322f
x_PM_DLLx1_ASAP7_75t_R%PD3 VSS N_MM9_s N_MM8_d N_PD3_1 PM_DLLx1_ASAP7_75t_R%PD3
cc_30 N_PD3_1 N_MM9_g 0.00772554f
cc_31 N_PD3_1 N_MM11_g 0.00775685f
x_PM_DLLx1_ASAP7_75t_R%PU1 VSS N_MM3_d N_MM1_s N_PU1_1 PM_DLLx1_ASAP7_75t_R%PU1
cc_32 N_PU1_1 N_MM3_g 0.0169868f
cc_33 N_PU1_1 N_MM1_g 0.0169686f
x_PM_DLLx1_ASAP7_75t_R%PD1 VSS N_MM5_d N_MM4_s N_PD1_5 N_PD1_4 N_PD1_1
+ PM_DLLx1_ASAP7_75t_R%PD1
cc_34 N_PD1_5 N_CLKN_2 0.000750294f
cc_35 N_PD1_5 N_MM10_g 0.0346381f
cc_36 N_PD1_4 N_D_1 0.000673808f
cc_37 N_PD1_4 N_D_4 0.000738828f
cc_38 N_PD1_4 N_MM3_g 0.0361067f
cc_39 N_PD1_5 N_CLKB_19 0.000497544f
cc_40 N_PD1_5 N_CLKB_1 0.00228924f
cc_41 N_PD1_5 N_MM1_g 0.0737342f
cc_42 N_PD1_1 N_MH_18 0.000162001f
cc_43 N_PD1_1 N_MH_6 0.00140674f
cc_44 N_PD1_1 N_MH_13 0.0031934f
x_PM_DLLx1_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_DLLx1_ASAP7_75t_R%noxref_18
cc_45 N_noxref_18_1 N_MM3_g 0.00135949f
cc_46 N_noxref_18_1 N_CLKB_18 0.000118156f
cc_47 N_noxref_18_1 N_CLKB_14 0.000701126f
cc_48 N_noxref_18_1 N_noxref_16_1 0.00769882f
cc_49 N_noxref_18_1 N_noxref_17_1 0.000465047f
x_PM_DLLx1_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_DLLx1_ASAP7_75t_R%noxref_19
cc_50 N_noxref_19_1 N_MM3_g 0.00136116f
cc_51 N_noxref_19_1 N_CLKB_18 0.000110294f
cc_52 N_noxref_19_1 N_CLKB_15 0.000665679f
cc_53 N_noxref_19_1 N_noxref_16_1 0.000465319f
cc_54 N_noxref_19_1 N_noxref_17_1 0.00769566f
cc_55 N_noxref_19_1 N_noxref_18_1 0.0012342f
x_PM_DLLx1_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_DLLx1_ASAP7_75t_R%noxref_16
cc_56 N_noxref_16_1 N_MM23_g 0.00394553f
cc_57 N_noxref_16_1 N_CLKB_4 0.000428447f
cc_58 N_noxref_16_1 N_CLKB_14 0.0270741f
x_PM_DLLx1_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_DLLx1_ASAP7_75t_R%noxref_17
cc_59 N_noxref_17_1 N_MM23_g 0.0040583f
cc_60 N_noxref_17_1 N_CLKB_5 0.000420714f
cc_61 N_noxref_17_1 N_CLKB_15 0.0270065f
cc_62 N_noxref_17_1 N_noxref_16_1 0.00141501f
x_PM_DLLx1_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_DLLx1_ASAP7_75t_R%noxref_21
cc_63 N_noxref_21_1 N_CLKB_6 0.00289337f
cc_64 N_noxref_21_1 N_NET085_11 0.0163862f
cc_65 N_noxref_21_1 N_MM7_g 0.00528057f
cc_66 N_noxref_21_1 N_noxref_20_1 0.00148265f
x_PM_DLLx1_ASAP7_75t_R%PD2 VSS N_MM10_s N_MM11_d N_PD2_4 N_PD2_5 N_PD2_1
+ PM_DLLx1_ASAP7_75t_R%PD2
cc_67 N_PD2_4 N_MM10_g 0.015171f
cc_68 N_PD2_5 N_CLKB_6 0.00128333f
cc_69 N_PD2_1 N_CLKB_2 0.00100177f
cc_70 N_PD2_1 N_MM9_g 0.00222097f
cc_71 N_PD2_4 N_MM9_g 0.00715002f
cc_72 N_PD2_5 N_MM9_g 0.0240095f
cc_73 N_PD2_5 N_MM11_g 0.0145993f
cc_74 N_PD2_1 N_MH_15 0.000609067f
cc_75 N_PD2_1 N_MH_20 0.00039116f
cc_76 N_PD2_1 N_MH_17 0.00041296f
cc_77 N_PD2_4 N_MH_5 0.000591818f
cc_78 N_PD2_1 N_MH_25 0.00211706f
x_PM_DLLx1_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_DLLx1_ASAP7_75t_R%noxref_23
cc_79 N_noxref_23_1 N_CLKB_6 0.000598937f
cc_80 N_noxref_23_1 N_MM25_g 0.00155737f
cc_81 N_noxref_23_1 N_noxref_20_1 0.00046945f
cc_82 N_noxref_23_1 N_noxref_21_1 0.00760944f
cc_83 N_noxref_23_1 N_noxref_22_1 0.0012286f
x_PM_DLLx1_ASAP7_75t_R%MH VSS N_MM7_g N_MM25_g N_MM4_d N_MM9_d N_MM1_d N_MM10_d
+ N_MH_21 N_MH_5 N_MH_16 N_MH_18 N_MH_15 N_MH_24 N_MH_26 N_MH_19 N_MH_20
+ N_MH_17 N_MH_6 N_MH_13 N_MH_14 N_MH_25 N_MH_1 N_MH_2 N_MH_22 N_MH_23
+ PM_DLLx1_ASAP7_75t_R%MH
cc_84 N_MH_21 N_MM10_g 0.000139334f
cc_85 N_MH_5 N_CLKN_21 0.000143656f
cc_86 N_MH_16 N_MM10_g 0.000177764f
cc_87 N_MH_18 N_CLKN_21 0.000235268f
cc_88 N_MH_15 N_MM10_g 0.0167259f
cc_89 N_MH_24 N_CLKN_21 0.00053907f
cc_90 N_MH_26 N_CLKN_27 0.000715688f
cc_91 N_MH_5 N_CLKN_2 0.000734988f
cc_92 N_MH_19 N_CLKN_21 0.000828006f
cc_93 N_MH_20 N_CLKN_21 0.00597797f
cc_94 N_MH_17 N_CLKN_27 0.000980364f
cc_95 N_MH_17 N_CLKN_21 0.00103345f
cc_96 N_MH_6 N_MM10_g 0.00110624f
cc_97 N_MH_5 N_MM10_g 0.00138094f
cc_98 N_MH_15 N_CLKN_2 0.00168951f
cc_99 N_MH_13 N_MM10_g 0.0535369f
cc_100 N_MH_13 N_CLKB_20 0.000112131f
cc_101 N_MH_17 N_CLKB_19 0.00134436f
cc_102 N_MH_16 N_MM1_g 0.000151732f
cc_103 N_MH_14 N_MM9_g 0.000170254f
cc_104 N_MH_5 N_CLKB_19 0.00152624f
cc_105 N_MH_19 N_CLKB_20 0.000242275f
cc_106 N_MH_15 N_MM1_g 0.0345508f
cc_107 N_MH_5 N_CLKB_1 0.000269762f
cc_108 N_MH_25 N_CLKB_20 0.000306266f
cc_109 N_MH_1 N_CLKB_6 0.00178862f
cc_110 N_MH_20 N_CLKB_23 0.000620396f
cc_111 N_MH_6 N_MM9_g 0.000632718f
cc_112 N_MH_26 N_CLKB_20 0.00070198f
cc_113 N_MH_21 N_CLKB_6 0.000717063f
cc_114 N_MH_15 N_CLKB_1 0.000794903f
cc_115 N_MH_20 N_CLKB_2 0.000887994f
cc_116 N_MH_5 N_MM1_g 0.00175046f
cc_117 N_MH_20 N_CLKB_20 0.00226127f
cc_118 N_MH_21 N_CLKB_20 0.00406011f
cc_119 N_MH_26 N_CLKB_23 0.00465639f
cc_120 N_MH_17 N_CLKB_23 0.00551743f
cc_121 N_MM7_g N_CLKB_6 0.00636423f
cc_122 N_MH_13 N_MM9_g 0.0370027f
cc_123 N_MH_18 N_MM11_g 7.28578e-20
cc_124 N_MH_2 N_MM11_g 8.57947e-20
cc_125 N_MH_13 N_MM11_g 0.000168215f
cc_126 N_MH_21 N_MM11_g 0.000180575f
cc_127 N_MM7_g N_NET085_3 0.000350173f
cc_128 N_MH_6 N_NET085_1 0.000445266f
cc_129 N_MH_26 N_NET085_16 0.00045396f
cc_130 N_MH_22 N_NET085_14 0.000493157f
cc_131 N_MH_21 N_NET085_13 0.000602008f
cc_132 N_MH_1 N_NET085_14 0.000742976f
cc_133 N_MH_21 N_NET085_1 0.000804847f
cc_134 N_MH_1 N_MM11_g 0.000911122f
cc_135 N_MH_23 N_NET085_15 0.000915448f
cc_136 N_MM7_g N_NET085_1 0.001082f
cc_137 N_MM7_g N_NET085_10 0.00660782f
cc_138 N_MM7_g N_NET085_11 0.00653853f
cc_139 N_MH_26 N_NET085_14 0.00260019f
cc_140 N_MH_21 N_NET085_12 0.00304766f
cc_141 N_MH_19 N_NET085_12 0.00360975f
cc_142 N_MH_21 N_NET085_14 0.00398201f
cc_143 N_MM7_g N_MM11_g 0.0293617f
x_PM_DLLx1_ASAP7_75t_R%CLK VSS CLK N_MM20_g N_CLK_8 N_CLK_6 N_CLK_1 N_CLK_7
+ N_CLK_5 N_CLK_4 PM_DLLx1_ASAP7_75t_R%CLK
x_PM_DLLx1_ASAP7_75t_R%D VSS D N_MM3_g N_D_4 N_D_5 N_D_6 N_D_1
+ PM_DLLx1_ASAP7_75t_R%D
cc_144 N_D_4 N_CLKN_21 0.000139517f
cc_145 N_D_4 N_CLKN_27 0.00279944f
x_PM_DLLx1_ASAP7_75t_R%NET085 VSS N_MM11_g N_MM6_d N_MM7_d N_NET085_16
+ N_NET085_11 N_NET085_1 N_NET085_4 N_NET085_14 N_NET085_3 N_NET085_13
+ N_NET085_15 N_NET085_10 N_NET085_12 PM_DLLx1_ASAP7_75t_R%NET085
cc_146 N_MM11_g N_CLKB_2 0.00015799f
cc_147 N_MM11_g N_CLKB_6 0.00516772f
cc_148 N_MM11_g N_CLKB_23 0.000190051f
cc_149 N_MM11_g N_CLKB_20 0.000253804f
cc_150 N_NET085_16 N_CLKB_6 0.000385253f
cc_151 N_NET085_11 N_CLKB_6 0.000386124f
cc_152 N_NET085_1 N_MM9_g 0.000414231f
cc_153 N_NET085_4 N_CLKB_6 0.000889986f
cc_154 N_NET085_14 N_CLKB_6 0.00128353f
cc_155 N_MM11_g N_MM9_g 0.0145065f
x_PM_DLLx1_ASAP7_75t_R%CLKN VSS N_MM23_g N_MM10_g N_MM20_d N_MM21_d N_CLKN_6
+ N_CLKN_5 N_CLKN_23 N_CLKN_13 N_CLKN_14 N_CLKN_1 N_CLKN_16 N_CLKN_18 N_CLKN_19
+ N_CLKN_17 N_CLKN_27 N_CLKN_25 N_CLKN_15 N_CLKN_21 N_CLKN_20 N_CLKN_26
+ N_CLKN_2 PM_DLLx1_ASAP7_75t_R%CLKN
cc_156 N_CLKN_6 N_MM20_g 0.00106627f
cc_157 N_CLKN_5 N_MM20_g 0.00109503f
cc_158 N_CLKN_23 N_MM20_g 0.000257621f
cc_159 N_CLKN_13 N_MM20_g 0.0112204f
cc_160 N_CLKN_14 N_MM20_g 0.0113266f
cc_161 N_CLKN_1 N_CLK_8 0.000419445f
cc_162 N_CLKN_16 N_CLK_8 0.000450651f
cc_163 N_CLKN_18 N_CLK_6 0.000686972f
cc_164 N_CLKN_23 N_CLK_1 0.000776704f
cc_165 N_CLKN_19 N_CLK_7 0.0015348f
cc_166 N_CLKN_17 N_CLK_5 0.00177807f
cc_167 N_CLKN_27 N_CLK_8 0.00202035f
cc_168 N_CLKN_23 N_CLK_8 0.00223928f
cc_169 N_CLKN_23 N_CLK_4 0.00230102f
cc_170 N_CLKN_25 N_CLK_6 0.0023102f
cc_171 N_CLKN_15 N_CLK_7 0.00242416f
cc_172 N_CLKN_1 N_CLK_1 0.0025247f
cc_173 N_CLKN_19 N_CLK_8 0.00264381f
cc_174 N_MM23_g N_MM20_g 0.0353315f
x_PM_DLLx1_ASAP7_75t_R%CLKB VSS N_MM1_g N_MM9_g N_MM23_d N_MM22_d N_CLKB_14
+ N_CLKB_5 N_CLKB_17 N_CLKB_4 N_CLKB_16 N_CLKB_21 N_CLKB_6 N_CLKB_15 N_CLKB_19
+ N_CLKB_18 N_CLKB_23 N_CLKB_2 N_CLKB_1 N_CLKB_22 N_CLKB_20
+ PM_DLLx1_ASAP7_75t_R%CLKB
cc_175 N_CLKB_14 N_CLK_5 8.44639e-20
cc_176 N_CLKB_5 N_CLK_5 0.00031786f
cc_177 N_CLKB_17 N_CLK_5 0.000160324f
cc_178 N_CLKB_4 N_CLK_5 0.000435192f
cc_179 N_CLKB_17 N_CLK_6 0.0010672f
cc_180 N_CLKB_16 N_CLK_5 0.00211738f
cc_181 N_CLKB_4 N_MM23_g 0.000858601f
cc_182 N_CLKB_21 N_MM23_g 0.000111867f
cc_183 N_CLKB_6 N_MM10_g 0.000169829f
cc_184 N_CLKB_15 N_MM23_g 0.0111469f
cc_185 N_CLKB_5 N_CLKN_25 0.000336745f
cc_186 N_CLKB_5 N_CLKN_1 0.00039569f
cc_187 N_CLKB_19 N_CLKN_27 0.000404678f
cc_188 N_CLKB_18 N_CLKN_20 0.00151691f
cc_189 N_CLKB_18 N_CLKN_19 0.000473746f
cc_190 N_CLKB_16 N_CLKN_26 0.000548968f
cc_191 N_CLKB_18 N_CLKN_27 0.000628391f
cc_192 N_CLKB_23 N_CLKN_21 0.000645472f
cc_193 N_CLKB_2 N_MM10_g 0.000669269f
cc_194 N_CLKB_1 N_CLKN_2 0.00215049f
cc_195 N_CLKB_15 N_CLKN_1 0.000897935f
cc_196 N_CLKB_5 N_MM23_g 0.00117264f
cc_197 N_MM1_g N_MM10_g 0.00162489f
cc_198 N_CLKB_18 N_CLKN_26 0.0041511f
cc_199 N_CLKB_19 N_CLKN_21 0.00457905f
cc_200 N_CLKB_17 N_CLKN_25 0.00559983f
cc_201 N_MM9_g N_MM10_g 0.00912894f
cc_202 N_CLKB_23 N_CLKN_27 0.0193279f
cc_203 N_CLKB_14 N_MM23_g 0.038949f
cc_204 N_CLKB_18 N_D_4 0.00352934f
cc_205 N_CLKB_21 N_D_5 0.000890482f
cc_206 N_CLKB_22 N_D_6 0.00089908f
cc_207 N_CLKB_23 N_D_6 0.000906642f
cc_208 N_CLKB_1 N_D_1 0.00273325f
cc_209 N_MM1_g N_MM3_g 0.00507026f
cc_210 N_CLKB_19 N_D_4 0.00920556f
*END of DLLx1_ASAP7_75t_R.pxi
.ENDS
** Design:	DLLx2_ASAP7_75t_R
* Created:	"Fri Aug 17 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "DLLx2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "DLLx2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_DLLx2_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00415905f
.ends

.subckt PM_DLLx2_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00424902f
.ends

.subckt PM_DLLx2_ASAP7_75t_R%PU1 VSS 2 4 1
c1 1 VSS 0.000968455f
r1 4 3 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3365 $Y2=0.2025
r2 2 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3195 $Y2=0.2025
r3 1 3 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3195 $Y=0.2025 $X2=0.3365 $Y2=0.2025
.ends

.subckt PM_DLLx2_ASAP7_75t_R%D VSS 9 3 4 5 6 1
c1 1 VSS 0.0065315f
c2 3 VSS 0.0833543f
c3 4 VSS 0.00563483f
c4 5 VSS 0.00674675f
c5 6 VSS 0.00728231f
r1 6 13 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.2340 $X2=0.2970 $Y2=0.2140
r2 12 13 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1735 $X2=0.2970 $Y2=0.2140
r3 11 12 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1735
r4 10 11 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1215 $X2=0.2970 $Y2=0.1350
r5 9 10 1.16595 $w=1.3e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1165 $X2=0.2970 $Y2=0.1215
r6 9 8 1.28254 $w=1.3e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1165 $X2=0.2970 $Y2=0.1110
r7 4 8 8.27824 $w=1.3e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0755 $X2=0.2970 $Y2=0.1110
r8 4 5 8.03069 $w=1.41392e-08 $l=3.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0755 $X2=0.2970 $Y2=0.0360
r9 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r10 1 11 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_DLLx2_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.0046906f
.ends

.subckt PM_DLLx2_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.041842f
.ends

.subckt PM_DLLx2_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.00467114f
.ends

.subckt PM_DLLx2_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.0417916f
.ends

.subckt PM_DLLx2_ASAP7_75t_R%PD3 VSS 2 4 1
c1 1 VSS 0.000929601f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0405 $X2=0.4905 $Y2=0.0405
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0405 $X2=0.4735 $Y2=0.0405
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4735 $Y=0.0405 $X2=0.4905 $Y2=0.0405
.ends

.subckt PM_DLLx2_ASAP7_75t_R%CLK VSS 11 3 8 6 1 4 7 5
c1 1 VSS 0.00252634f
c2 3 VSS 0.0597163f
c3 4 VSS 0.000784621f
c4 5 VSS 0.00424231f
c5 6 VSS 0.00413935f
c6 7 VSS 0.00189552f
c7 8 VSS 0.00176723f
r1 6 17 2.40741 $w=2.45e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.1980 $X2=0.1080 $Y2=0.1710
r2 5 15 4.50612 $w=2.06667e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0630 $X2=0.1080 $Y2=0.0990
r3 16 17 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.1710 $X2=0.1080 $Y2=0.1710
r4 8 13 1.35805 $w=2.83333e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1710 $X2=0.0810 $Y2=0.1485
r5 8 16 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1710 $X2=0.0945 $Y2=0.1710
r6 14 15 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.0990 $X2=0.1080 $Y2=0.0990
r7 7 10 0.483592 $w=3.42308e-08 $l=1.87e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0990 $X2=0.0810 $Y2=0.1177
r8 7 14 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0990 $X2=0.0945 $Y2=0.0990
r9 11 12 0.874462 $w=1.3e-08 $l=3.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1227
r10 11 10 0.291487 $w=1.3e-08 $l=1.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1177
r11 4 12 2.85657 $w=1.3e-08 $l=1.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1227
r12 4 13 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1485
r13 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r14 1 4 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_DLLx2_ASAP7_75t_R%PD1 VSS 7 10 5 4 1
c1 1 VSS 0.00934545f
c2 4 VSS 0.00316938f
c3 5 VSS 0.00186596f
r1 10 9 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r2 8 9 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r3 5 8 0.123457 $w=8.1e-08 $l=1e-08 $layer=N_src_drn $thickness=1e-09 $X=0.3780
+ $Y=0.0675 $X2=0.3880 $Y2=0.0675
r4 4 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3220 $Y2=0.0675
r5 7 4 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r6 1 5 1e-05
.ends

.subckt PM_DLLx2_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.00385186f
.ends

.subckt PM_DLLx2_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.00302765f
.ends

.subckt PM_DLLx2_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.00457728f
.ends

.subckt PM_DLLx2_ASAP7_75t_R%PD2 VSS 7 13 4 5 1
c1 1 VSS 0.00713406f
c2 4 VSS 0.00187814f
c3 5 VSS 0.00233943f
r1 13 12 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r2 5 12 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4880 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r3 10 5 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4725
+ $Y=0.2295 $X2=0.4860 $Y2=0.2295
r4 9 10 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4590
+ $Y=0.2295 $X2=0.4725 $Y2=0.2295
r5 8 9 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4455
+ $Y=0.2295 $X2=0.4590 $Y2=0.2295
r6 1 8 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4320
+ $Y=0.2295 $X2=0.4455 $Y2=0.2295
r7 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2295 $X2=0.4300 $Y2=0.2295
r8 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2295 $X2=0.4175 $Y2=0.2295
.ends

.subckt PM_DLLx2_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.00487759f
.ends

.subckt PM_DLLx2_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.00511776f
.ends

.subckt PM_DLLx2_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.00488042f
.ends

.subckt PM_DLLx2_ASAP7_75t_R%NET085 VSS 9 35 40 4 16 11 1 14 10 3 13 15 12 17
c1 1 VSS 0.00286915f
c2 3 VSS 0.00565906f
c3 4 VSS 0.00633095f
c4 9 VSS 0.0374877f
c5 10 VSS 0.00324794f
c6 11 VSS 0.00343435f
c7 12 VSS 0.00127673f
c8 13 VSS 0.00859887f
c9 14 VSS 0.00297262f
c10 15 VSS 0.00281155f
c11 16 VSS 0.00574037f
c12 17 VSS 0.00269091f
r1 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2295 $X2=0.5920 $Y2=0.2295
r2 40 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.2295 $X2=0.5795 $Y2=0.2295
r3 4 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2295
+ $X2=0.5940 $Y2=0.2340
r4 37 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.2340 $X2=0.6075 $Y2=0.2340
r5 16 33 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.2340 $X2=0.6210 $Y2=0.2140
r6 16 38 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.2340 $X2=0.6075 $Y2=0.2340
r7 10 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.0405 $X2=0.5920 $Y2=0.0405
r8 35 10 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0405 $X2=0.5795 $Y2=0.0405
r9 32 33 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1850 $X2=0.6210 $Y2=0.2140
r10 31 32 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1660 $X2=0.6210 $Y2=0.1850
r11 30 31 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1525 $X2=0.6210 $Y2=0.1660
r12 29 30 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1310 $X2=0.6210 $Y2=0.1525
r13 28 29 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1095 $X2=0.6210 $Y2=0.1310
r14 27 28 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0935 $X2=0.6210 $Y2=0.1095
r15 14 17 5.69636 $w=1.58e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.0675 $X2=0.6210 $Y2=0.0360
r16 14 27 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0675 $X2=0.6210 $Y2=0.0935
r17 3 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0405
+ $X2=0.5940 $Y2=0.0360
r18 17 26 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.0360 $X2=0.6075 $Y2=0.0360
r19 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0360 $X2=0.6075 $Y2=0.0360
r20 24 25 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5825
+ $Y=0.0360 $X2=0.5940 $Y2=0.0360
r21 13 15 7.2121 $w=1.41842e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5510 $Y=0.0360 $X2=0.5130 $Y2=0.0360
r22 13 24 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5510
+ $Y=0.0360 $X2=0.5825 $Y2=0.0360
r23 12 22 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0590 $X2=0.5130 $Y2=0.0820
r24 12 15 3.71425 $w=1.68348e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.0590 $X2=0.5130 $Y2=0.0360
r25 1 19 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.5130
+ $Y=0.0820 $X2=0.5130 $Y2=0.0820
r26 1 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.0820
+ $X2=0.5130 $Y2=0.0820
r27 9 19 0.314665 $w=2.27e-07 $l=5.3e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5130 $Y2=0.0820
.ends

.subckt PM_DLLx2_ASAP7_75t_R%Q VSS 35 23 38 51 53 1 18 17 2 13 16 14 15 19 4 3
c1 1 VSS 0.00841373f
c2 2 VSS 0.00853601f
c3 3 VSS 0.00756745f
c4 4 VSS 0.00763753f
c5 13 VSS 0.00348946f
c6 14 VSS 0.00347753f
c7 15 VSS 0.00403083f
c8 16 VSS 0.00347266f
c9 17 VSS 0.0137612f
c10 18 VSS 0.0139032f
c11 19 VSS 0.0030425f
c12 20 VSS 0.00270003f
c13 21 VSS 0.00273657f
r1 53 52 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.2025 $X2=0.7165 $Y2=0.2025
r2 15 52 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7040 $Y=0.2025 $X2=0.7165 $Y2=0.2025
r3 16 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.2025 $X2=0.8080 $Y2=0.2025
r4 51 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.2025 $X2=0.7955 $Y2=0.2025
r5 2 43 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7020 $Y=0.2295
+ $X2=0.7020 $Y2=0.2340
r6 4 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8100 $Y=0.2025
+ $X2=0.8100 $Y2=0.2340
r7 43 44 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.2340 $X2=0.7425 $Y2=0.2340
r8 41 44 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.2340 $X2=0.7425 $Y2=0.2340
r9 39 40 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.2340 $X2=0.8240 $Y2=0.2340
r10 18 39 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7965
+ $Y=0.2340 $X2=0.8100 $Y2=0.2340
r11 18 41 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7965
+ $Y=0.2340 $X2=0.7830 $Y2=0.2340
r12 21 36 0.624487 $w=2.20462e-08 $l=9.8e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.8380 $Y=0.2340 $X2=0.8380 $Y2=0.2242
r13 21 40 1.61554 $w=1.62143e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8380 $Y=0.2340 $X2=0.8240 $Y2=0.2340
r14 14 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.0675 $X2=0.8080 $Y2=0.0675
r15 38 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.0675 $X2=0.7955 $Y2=0.0675
r16 35 36 0.291487 $w=1.3e-08 $l=1.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.8380
+ $Y=0.2230 $X2=0.8380 $Y2=0.2242
r17 35 34 6.58761 $w=1.3e-08 $l=2.83e-08 $layer=M1 $thickness=3.6e-08 $X=0.8380
+ $Y=0.2230 $X2=0.8380 $Y2=0.1947
r18 33 34 15.4488 $w=1.3e-08 $l=6.62e-08 $layer=M1 $thickness=3.6e-08 $X=0.8380
+ $Y=0.1285 $X2=0.8380 $Y2=0.1947
r19 19 20 5.69636 $w=1.58e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8380 $Y=0.0675 $X2=0.8380 $Y2=0.0360
r20 19 33 14.2246 $w=1.3e-08 $l=6.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.8380
+ $Y=0.0675 $X2=0.8380 $Y2=0.1285
r21 3 31 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8100 $Y=0.0675
+ $X2=0.8100 $Y2=0.0360
r22 20 32 1.61554 $w=1.62143e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8380 $Y=0.0360 $X2=0.8240 $Y2=0.0360
r23 31 32 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.8100
+ $Y=0.0360 $X2=0.8240 $Y2=0.0360
r24 30 31 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7965
+ $Y=0.0360 $X2=0.8100 $Y2=0.0360
r25 29 30 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.0360 $X2=0.7965 $Y2=0.0360
r26 28 29 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.7425
+ $Y=0.0360 $X2=0.7830 $Y2=0.0360
r27 27 28 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.0360 $X2=0.7425 $Y2=0.0360
r28 17 27 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6905
+ $Y=0.0360 $X2=0.7020 $Y2=0.0360
r29 13 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7020 $Y=0.0405
+ $X2=0.7020 $Y2=0.0360
r30 1 13 12.9669 $w=2.02e-08 $l=2.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.7020 $Y=0.0625 $X2=0.7020 $Y2=0.0405
r31 23 22 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.0675 $X2=0.7165 $Y2=0.0675
r32 13 22 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7040 $Y=0.0675 $X2=0.7165 $Y2=0.0675
r33 2 15 1e-05
.ends

.subckt PM_DLLx2_ASAP7_75t_R%CLKN VSS 11 12 66 68 6 5 23 13 14 1 16 18 19 17 27
+ 25 15 21 20 26 2
c1 1 VSS 0.00166015f
c2 2 VSS 7.18467e-20
c3 5 VSS 0.00755214f
c4 6 VSS 0.00759316f
c5 11 VSS 0.0597516f
c6 12 VSS 0.00453873f
c7 13 VSS 0.00561806f
c8 14 VSS 0.00562522f
c9 15 VSS 0.0048817f
c10 16 VSS 0.00316121f
c11 17 VSS 0.00479583f
c12 18 VSS 0.00459222f
c13 19 VSS 0.000422747f
c14 20 VSS 0.000372814f
c15 21 VSS 0.000774523f
c16 22 VSS 0.00358581f
c17 23 VSS 0.00143173f
c18 24 VSS 0.00361511f
c19 25 VSS 0.000791544f
c20 26 VSS 0.00040304f
c21 27 VSS 0.0135925f
r1 68 67 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r2 14 67 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r3 66 65 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r4 13 65 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r5 6 63 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0550 $Y2=0.2340
r6 5 60 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0550 $Y2=0.0360
r7 62 63 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.2340 $X2=0.0550 $Y2=0.2340
r8 18 62 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0460 $Y2=0.2340
r9 18 24 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0180 $Y2=0.2340
r10 59 60 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.0360 $X2=0.0550 $Y2=0.0360
r11 17 59 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0460 $Y2=0.0360
r12 17 22 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0180 $Y2=0.0360
r13 12 57 5.63117 $w=1.26721e-07 $l=2e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4050 $Y2=0.1330
r14 24 56 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.2340 $X2=0.0180 $Y2=0.2070
r15 22 55 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.0360 $X2=0.0180 $Y2=0.0630
r16 2 57 6.49795 $w=1.53e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08 $X=0.4050
+ $Y=0.1440 $X2=0.4050 $Y2=0.1330
r17 16 23 3.9134 $w=1.47857e-08 $l=2.25499e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1755 $X2=0.0165 $Y2=0.1530
r18 16 56 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1755 $X2=0.0180 $Y2=0.2070
r19 54 55 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0990 $X2=0.0180 $Y2=0.0630
r20 15 23 3.9134 $w=1.47857e-08 $l=2.25499e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1305 $X2=0.0165 $Y2=0.1530
r21 15 54 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1305 $X2=0.0180 $Y2=0.0990
r22 52 57 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1440
+ $X2=0.4050 $Y2=0.1330
r23 21 52 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1160 $X2=0.4050 $Y2=0.1440
r24 49 50 1.90199 $w=1.38333e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.0255 $Y=0.1530 $X2=0.0345 $Y2=0.1530
r25 23 49 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0165
+ $Y=0.1530 $X2=0.0255 $Y2=0.1530
r26 25 41 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1980 $X2=0.1890 $Y2=0.1755
r27 47 52 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4050 $Y=0.1530
+ $X2=0.4050 $Y2=0.1440
r28 46 47 21.5701 $w=1.3e-08 $l=9.25e-08 $layer=M2 $thickness=3.6e-08 $X=0.3125
+ $Y=0.1530 $X2=0.4050 $Y2=0.1530
r29 45 46 23.0858 $w=1.3e-08 $l=9.9e-08 $layer=M2 $thickness=3.6e-08 $X=0.2135
+ $Y=0.1530 $X2=0.3125 $Y2=0.1530
r30 44 45 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1530 $X2=0.2135 $Y2=0.1530
r31 43 44 18.1888 $w=1.3e-08 $l=7.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.1110
+ $Y=0.1530 $X2=0.1890 $Y2=0.1530
r32 42 43 18.1888 $w=1.3e-08 $l=7.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.0330
+ $Y=0.1530 $X2=0.1110 $Y2=0.1530
r33 42 50 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.0330 $Y=0.1530
+ $X2=0.0345 $Y2=0.1530
r34 27 42 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.0215
+ $Y=0.1530 $X2=0.0330 $Y2=0.1530
r35 40 41 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1575 $X2=0.1890 $Y2=0.1755
r36 20 26 1.49895 $w=1.95333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1485 $X2=0.1890 $Y2=0.1350
r37 20 40 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1485 $X2=0.1890 $Y2=0.1575
r38 20 44 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1890 $Y=0.1485
+ $X2=0.1890 $Y2=0.1530
r39 26 39 2.6649 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1705 $Y2=0.1350
r40 38 39 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.1545
+ $Y=0.1350 $X2=0.1705 $Y2=0.1350
r41 37 38 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1455
+ $Y=0.1350 $X2=0.1545 $Y2=0.1350
r42 19 37 1.16595 $w=1.3e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1405
+ $Y=0.1350 $X2=0.1455 $Y2=0.1350
r43 35 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1555 $Y=0.1350
+ $X2=0.1545 $Y2=0.1350
r44 34 35 4.72579 $w=1.53e-08 $l=8e-09 $layer=LIG $thickness=4.8e-08 $X=0.1475
+ $Y=0.1350 $X2=0.1555 $Y2=0.1350
r45 32 34 1.73797 $w=1.72143e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1440 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r46 1 32 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.1340
+ $Y=0.1350 $X2=0.1440 $Y2=0.1350
r47 11 1 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1340 $Y2=0.1350
r48 11 34 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r49 6 14 1e-05
r50 5 13 1e-05
.ends

.subckt PM_DLLx2_ASAP7_75t_R%CLKB VSS 12 13 71 73 14 5 17 4 16 21 6 15 19 18 23
+ 2 1 22 20
c1 1 VSS 0.000282427f
c2 2 VSS 9.10164e-20
c3 4 VSS 0.00691117f
c4 5 VSS 0.00721883f
c5 6 VSS 0.00500393f
c6 12 VSS 0.00528809f
c7 13 VSS 0.00505164f
c8 14 VSS 0.00642769f
c9 15 VSS 0.00638157f
c10 16 VSS 0.0100164f
c11 17 VSS 0.00897636f
c12 18 VSS 0.00623091f
c13 19 VSS 0.00120388f
c14 20 VSS 0.00152188f
c15 21 VSS 0.0031578f
c16 22 VSS 0.00304667f
c17 23 VSS 0.0111991f
r1 15 5 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1600 $Y2=0.2160
r2 73 15 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r3 14 4 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1600 $Y2=0.0540
r4 71 14 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r5 5 66 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r6 4 63 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r7 2 54 5.67512 $w=2.4e-08 $l=5e-09 $layer=LISD $thickness=4.02632e-08
+ $X=0.4590 $Y=0.1790 $X2=0.4640 $Y2=0.1790
r8 13 2 2.88446 $w=1.16273e-07 $l=4.4e-08 $layer=LIG $thickness=5.16364e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4590 $Y2=0.1790
r9 66 67 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1845 $Y2=0.2340
r10 17 22 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.2340 $X2=0.2430 $Y2=0.2340
r11 17 67 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.1845 $Y2=0.2340
r12 63 64 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1845 $Y2=0.0360
r13 16 21 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.0360 $X2=0.2430 $Y2=0.0360
r14 16 64 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.1845 $Y2=0.0360
r15 52 54 11.0623 $w=2.14976e-08 $l=2.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4845 $Y=0.1790 $X2=0.4640 $Y2=0.1790
r16 51 52 8.84105 $w=2.02e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4995 $Y=0.1790 $X2=0.4845 $Y2=0.1790
r17 6 49 6.18874 $w=2.02e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5025 $Y=0.1790 $X2=0.5130 $Y2=0.1790
r18 6 51 1.76821 $w=2.02e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.5025
+ $Y=0.1790 $X2=0.4995 $Y2=0.1790
r19 22 46 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2430 $Y2=0.2160
r20 21 43 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0360 $X2=0.2430 $Y2=0.0630
r21 47 49 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5130 $Y=0.1845
+ $X2=0.5130 $Y2=0.1790
r22 20 47 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1680 $X2=0.5130 $Y2=0.1845
r23 45 46 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2025 $X2=0.2430 $Y2=0.2160
r24 44 45 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1935 $X2=0.2430 $Y2=0.2025
r25 42 43 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0990 $X2=0.2430 $Y2=0.0630
r26 41 42 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1215 $X2=0.2430 $Y2=0.0990
r27 40 44 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1845 $X2=0.2430 $Y2=0.1935
r28 18 40 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1530 $X2=0.2430 $Y2=0.1845
r29 18 41 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1530 $X2=0.2430 $Y2=0.1215
r30 38 47 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.5130 $Y=0.1890
+ $X2=0.5130 $Y2=0.1845
r31 37 38 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.4770
+ $Y=0.1890 $X2=0.5130 $Y2=0.1890
r32 36 37 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M2 $thickness=3.6e-08 $X=0.4320
+ $Y=0.1890 $X2=0.4770 $Y2=0.1890
r33 35 36 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M2 $thickness=3.6e-08 $X=0.3870
+ $Y=0.1890 $X2=0.4320 $Y2=0.1890
r34 34 35 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1890 $X2=0.3870 $Y2=0.1890
r35 33 34 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1890 $X2=0.3510 $Y2=0.1890
r36 32 33 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1890 $X2=0.2970 $Y2=0.1890
r37 32 40 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.2430 $Y=0.1890
+ $X2=0.2430 $Y2=0.1845
r38 23 32 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.2315
+ $Y=0.1890 $X2=0.2430 $Y2=0.1890
r39 29 34 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.3510 $Y=0.1890
+ $X2=0.3510 $Y2=0.1890
r40 28 29 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1620 $X2=0.3510 $Y2=0.1890
r41 27 28 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1620
r42 19 27 4.4306 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1160 $X2=0.3510 $Y2=0.1350
r43 12 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r44 1 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
.ends

.subckt PM_DLLx2_ASAP7_75t_R%MH VSS 11 12 13 72 76 81 85 22 5 17 19 16 25 27 20
+ 21 18 6 14 15 26 1 23 2 24
c1 1 VSS 0.000312313f
c2 2 VSS 0.00932051f
c3 5 VSS 0.00620842f
c4 6 VSS 0.00504477f
c5 11 VSS 0.0368722f
c6 12 VSS 0.080066f
c7 13 VSS 0.0801317f
c8 14 VSS 0.00410542f
c9 15 VSS 0.000930242f
c10 16 VSS 0.00452723f
c11 17 VSS 0.00092506f
c12 18 VSS 0.00790275f
c13 19 VSS 0.0039096f
c14 20 VSS 0.00122945f
c15 21 VSS 0.000699644f
c16 22 VSS 0.000513074f
c17 23 VSS 0.00284023f
c18 24 VSS 0.00250965f
c19 25 VSS 5.91466e-20
c20 26 VSS 0.00245709f
c21 27 VSS 0.0123703f
r1 85 84 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r2 83 84 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r3 16 83 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3760 $Y=0.2295 $X2=0.3880 $Y2=0.2295
r4 17 16 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2295 $X2=0.3760 $Y2=0.2295
r5 79 80 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r6 81 79 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.1890 $X2=0.3635 $Y2=0.1890
r7 16 80 0.185185 $w=5.4e-08 $l=1e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r8 12 65 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=0.7290
+ $Y=0.1350 $X2=0.7290 $Y2=0.1360
r9 13 58 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.7830 $Y=0.1350 $X2=0.7830 $Y2=0.1360
r10 76 75 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r11 74 75 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4420 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r12 6 74 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4300 $Y=0.0405 $X2=0.4420 $Y2=0.0405
r13 15 6 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0405 $X2=0.4300 $Y2=0.0405
r14 14 6 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0810 $X2=0.4300 $Y2=0.0810
r15 72 14 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0810 $X2=0.4175 $Y2=0.0810
r16 68 16 15.0298 $w=2.02e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.3780 $Y=0.2045 $X2=0.3780 $Y2=0.1790
r17 5 53 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2295
+ $X2=0.3780 $Y2=0.2340
r18 5 68 14.7351 $w=2.02e-08 $l=2.5e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.3780 $Y=0.2295 $X2=0.3780 $Y2=0.2045
r19 63 65 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7415 $Y=0.1360 $X2=0.7290 $Y2=0.1360
r20 62 63 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7560 $Y=0.1360 $X2=0.7415 $Y2=0.1360
r21 60 62 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7705 $Y=0.1360 $X2=0.7560 $Y2=0.1360
r22 2 58 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.7735
+ $Y=0.1360 $X2=0.7830 $Y2=0.1360
r23 2 60 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.7735 $Y=0.1360 $X2=0.7705 $Y2=0.1360
r24 6 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0405
+ $X2=0.4320 $Y2=0.0360
r25 53 54 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r26 51 54 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r27 18 26 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4320 $Y=0.2340 $X2=0.4590 $Y2=0.2340
r28 18 51 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4050 $Y2=0.2340
r29 49 58 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7830 $Y=0.1445
+ $X2=0.7830 $Y2=0.1360
r30 23 49 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1085 $X2=0.7830 $Y2=0.1445
r31 19 24 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4320 $Y=0.0360 $X2=0.4590 $Y2=0.0360
r32 26 44 3.01468 $w=1.741e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4590 $Y2=0.2140
r33 47 49 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.7830 $Y=0.1530
+ $X2=0.7830 $Y2=0.1445
r34 46 47 30.8976 $w=1.3e-08 $l=1.325e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.6505 $Y=0.1530 $X2=0.7830 $Y2=0.1530
r35 45 46 35.678 $w=1.3e-08 $l=1.53e-07 $layer=M2 $thickness=3.6e-08 $X=0.4975
+ $Y=0.1530 $X2=0.6505 $Y2=0.1530
r36 27 45 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M2 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1530 $X2=0.4975 $Y2=0.1530
r37 27 40 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4590 $Y=0.1530
+ $X2=0.4590 $Y2=0.1530
r38 24 39 6.51253 $w=1.552e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4590 $Y2=0.0710
r39 43 44 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2015 $X2=0.4590 $Y2=0.2140
r40 42 43 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1825 $X2=0.4590 $Y2=0.2015
r41 41 42 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1635 $X2=0.4590 $Y2=0.1825
r42 40 41 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1530 $X2=0.4590 $Y2=0.1635
r43 21 40 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1420 $X2=0.4590 $Y2=0.1530
r44 21 25 1.38478 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1420 $X2=0.4590 $Y2=0.1310
r45 38 39 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1015 $X2=0.4590 $Y2=0.0710
r46 20 25 2.78392 $w=1.56471e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1140 $X2=0.4590 $Y2=0.1310
r47 20 38 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1140 $X2=0.4590 $Y2=0.1015
r48 25 37 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1310 $X2=0.4860 $Y2=0.1310
r49 36 37 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1310 $X2=0.4860 $Y2=0.1310
r50 22 34 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.5395
+ $Y=0.1310 $X2=0.5660 $Y2=0.1310
r51 22 36 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.5395
+ $Y=0.1310 $X2=0.5130 $Y2=0.1310
r52 1 31 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.5670
+ $Y=0.1310 $X2=0.5670 $Y2=0.1310
r53 1 34 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1310
+ $X2=0.5660 $Y2=0.1310
r54 11 31 0.314665 $w=2.27e-07 $l=4e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5670 $Y=0.1350 $X2=0.5670 $Y2=0.1310
.ends


*
.SUBCKT DLLx2_ASAP7_75t_R VSS VDD CLK D Q
*
* VSS VSS
* VDD VDD
* CLK CLK
* D D
* Q Q
*
*

MM20 N_MM20_d N_MM20_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM23 N_MM23_d N_MM22_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM10_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM6 N_MM6_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM24 N_MM24_d N_MM25_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@2 N_MM24@2_d N_MM25@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM21 N_MM21_d N_MM20_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM22 N_MM22_d N_MM22_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM25 N_MM25_d N_MM25_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@2 N_MM25@2_d N_MM25@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "DLLx2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "DLLx2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_DLLx2_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_DLLx2_ASAP7_75t_R%noxref_15
cc_1 N_noxref_15_1 N_MM20_g 0.00366574f
cc_2 N_noxref_15_1 N_CLKN_16 0.000199342f
cc_3 N_noxref_15_1 N_CLKN_6 0.000504268f
cc_4 N_noxref_15_1 N_CLKN_14 0.0280996f
cc_5 N_noxref_15_1 N_noxref_14_1 0.00204873f
x_PM_DLLx2_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_DLLx2_ASAP7_75t_R%noxref_14
cc_6 N_noxref_14_1 N_MM20_g 0.00368079f
cc_7 N_noxref_14_1 N_CLKN_15 0.000315662f
cc_8 N_noxref_14_1 N_CLKN_5 0.000503546f
cc_9 N_noxref_14_1 N_CLKN_13 0.0279133f
x_PM_DLLx2_ASAP7_75t_R%PU1 VSS N_MM3_d N_MM1_s N_PU1_1 PM_DLLx2_ASAP7_75t_R%PU1
cc_10 N_PU1_1 N_MM3_g 0.0169893f
cc_11 N_PU1_1 N_MM1_g 0.0169659f
x_PM_DLLx2_ASAP7_75t_R%D VSS D N_MM3_g N_D_4 N_D_5 N_D_6 N_D_1
+ PM_DLLx2_ASAP7_75t_R%D
cc_12 N_D_4 N_CLKN_21 0.000245177f
cc_13 N_D_4 N_CLKN_27 0.00269342f
x_PM_DLLx2_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_DLLx2_ASAP7_75t_R%noxref_16
cc_14 N_noxref_16_1 N_MM22_g 0.00394553f
cc_15 N_noxref_16_1 N_CLKB_4 0.000428447f
cc_16 N_noxref_16_1 N_CLKB_14 0.0270742f
x_PM_DLLx2_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_DLLx2_ASAP7_75t_R%noxref_19
cc_17 N_noxref_19_1 N_MM3_g 0.00136116f
cc_18 N_noxref_19_1 N_CLKB_18 0.000110505f
cc_19 N_noxref_19_1 N_CLKB_15 0.000665197f
cc_20 N_noxref_19_1 N_noxref_16_1 0.00046532f
cc_21 N_noxref_19_1 N_noxref_17_1 0.00769567f
cc_22 N_noxref_19_1 N_noxref_18_1 0.00123419f
x_PM_DLLx2_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_DLLx2_ASAP7_75t_R%noxref_17
cc_23 N_noxref_17_1 N_CLKN_1 0.000395326f
cc_24 N_noxref_17_1 N_MM22_g 0.00366298f
cc_25 N_noxref_17_1 N_CLKB_5 0.000420714f
cc_26 N_noxref_17_1 N_CLKB_15 0.0270062f
cc_27 N_noxref_17_1 N_noxref_16_1 0.00141501f
x_PM_DLLx2_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_DLLx2_ASAP7_75t_R%noxref_18
cc_28 N_noxref_18_1 N_MM3_g 0.00135947f
cc_29 N_noxref_18_1 N_CLKB_18 0.000116624f
cc_30 N_noxref_18_1 N_CLKB_14 0.000701358f
cc_31 N_noxref_18_1 N_noxref_16_1 0.00769878f
cc_32 N_noxref_18_1 N_noxref_17_1 0.000465046f
x_PM_DLLx2_ASAP7_75t_R%PD3 VSS N_MM9_s N_MM8_d N_PD3_1 PM_DLLx2_ASAP7_75t_R%PD3
cc_33 N_PD3_1 N_MM9_g 0.00772678f
cc_34 N_PD3_1 N_MM11_g 0.00775685f
x_PM_DLLx2_ASAP7_75t_R%CLK VSS CLK N_MM20_g N_CLK_8 N_CLK_6 N_CLK_1 N_CLK_4
+ N_CLK_7 N_CLK_5 PM_DLLx2_ASAP7_75t_R%CLK
x_PM_DLLx2_ASAP7_75t_R%PD1 VSS N_MM5_d N_MM4_s N_PD1_5 N_PD1_4 N_PD1_1
+ PM_DLLx2_ASAP7_75t_R%PD1
cc_35 N_PD1_5 N_CLKN_2 0.000750248f
cc_36 N_PD1_5 N_MM10_g 0.0346358f
cc_37 N_PD1_4 N_D_1 0.000673767f
cc_38 N_PD1_4 N_D_4 0.00073878f
cc_39 N_PD1_4 N_MM3_g 0.0361045f
cc_40 N_PD1_5 N_CLKB_19 0.000497517f
cc_41 N_PD1_5 N_CLKB_1 0.0022891f
cc_42 N_PD1_5 N_MM1_g 0.0737372f
cc_43 N_PD1_1 N_MH_19 0.000161991f
cc_44 N_PD1_1 N_MH_6 0.00140665f
cc_45 N_PD1_1 N_MH_14 0.0031962f
x_PM_DLLx2_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_DLLx2_ASAP7_75t_R%noxref_20
cc_46 N_noxref_20_1 N_NET085_10 0.0170268f
cc_47 N_noxref_20_1 N_MM7_g 0.00582769f
cc_48 N_noxref_20_1 N_Q_13 0.000778394f
x_PM_DLLx2_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_DLLx2_ASAP7_75t_R%noxref_21
cc_49 N_noxref_21_1 N_CLKB_6 0.00289368f
cc_50 N_noxref_21_1 N_NET085_11 0.0163748f
cc_51 N_noxref_21_1 N_MM7_g 0.00528337f
cc_52 N_noxref_21_1 N_Q_15 0.000595359f
cc_53 N_noxref_21_1 N_noxref_20_1 0.00148436f
x_PM_DLLx2_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_DLLx2_ASAP7_75t_R%noxref_22
cc_54 N_noxref_22_1 N_NET085_10 0.00057322f
cc_55 N_noxref_22_1 N_MM25_g 0.00156965f
cc_56 N_noxref_22_1 N_Q_13 0.0372726f
cc_57 N_noxref_22_1 N_noxref_20_1 0.00775661f
cc_58 N_noxref_22_1 N_noxref_21_1 0.000455535f
x_PM_DLLx2_ASAP7_75t_R%PD2 VSS N_MM10_s N_MM11_d N_PD2_4 N_PD2_5 N_PD2_1
+ PM_DLLx2_ASAP7_75t_R%PD2
cc_59 N_PD2_4 N_MM10_g 0.0151666f
cc_60 N_PD2_5 N_CLKB_6 0.00128291f
cc_61 N_PD2_1 N_CLKB_2 0.00100148f
cc_62 N_PD2_1 N_MM9_g 0.00222032f
cc_63 N_PD2_4 N_MM9_g 0.00714792f
cc_64 N_PD2_5 N_MM9_g 0.0240218f
cc_65 N_PD2_5 N_MM11_g 0.014595f
cc_66 N_PD2_1 N_MH_16 0.000608888f
cc_67 N_PD2_1 N_MH_21 0.000391045f
cc_68 N_PD2_1 N_MH_18 0.000412839f
cc_69 N_PD2_4 N_MH_5 0.000591645f
cc_70 N_PD2_1 N_MH_26 0.00212147f
x_PM_DLLx2_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_DLLx2_ASAP7_75t_R%noxref_23
cc_71 N_noxref_23_1 N_CLKB_6 0.000597063f
cc_72 N_noxref_23_1 N_MM25_g 0.00150742f
cc_73 N_noxref_23_1 N_Q_15 0.0371896f
cc_74 N_noxref_23_1 N_noxref_20_1 0.000465679f
cc_75 N_noxref_23_1 N_noxref_21_1 0.00760048f
cc_76 N_noxref_23_1 N_noxref_22_1 0.00123903f
x_PM_DLLx2_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_DLLx2_ASAP7_75t_R%noxref_24
cc_77 N_noxref_24_1 N_MM25@2_g 0.00151672f
cc_78 N_noxref_24_1 N_Q_3 0.0005012f
cc_79 N_noxref_24_1 N_Q_14 0.0374856f
x_PM_DLLx2_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_DLLx2_ASAP7_75t_R%noxref_25
cc_80 N_noxref_25_1 N_MM25@2_g 0.00153281f
cc_81 N_noxref_25_1 N_Q_4 0.000501839f
cc_82 N_noxref_25_1 N_Q_16 0.0377627f
cc_83 N_noxref_25_1 N_noxref_24_1 0.00176462f
x_PM_DLLx2_ASAP7_75t_R%NET085 VSS N_MM11_g N_MM6_d N_MM7_d N_NET085_4
+ N_NET085_16 N_NET085_11 N_NET085_1 N_NET085_14 N_NET085_10 N_NET085_3
+ N_NET085_13 N_NET085_15 N_NET085_12 N_NET085_17 PM_DLLx2_ASAP7_75t_R%NET085
cc_84 N_MM11_g N_CLKB_2 0.00015799f
cc_85 N_MM11_g N_CLKB_6 0.00486101f
cc_86 N_MM11_g N_CLKB_23 0.00018317f
cc_87 N_MM11_g N_CLKB_20 0.000253804f
cc_88 N_NET085_4 N_CLKB_6 0.00119662f
cc_89 N_NET085_16 N_CLKB_6 0.000372952f
cc_90 N_NET085_11 N_CLKB_6 0.000379122f
cc_91 N_NET085_1 N_MM9_g 0.000414231f
cc_92 N_NET085_14 N_CLKB_6 0.00128164f
cc_93 N_MM11_g N_MM9_g 0.0144986f
x_PM_DLLx2_ASAP7_75t_R%Q VSS Q N_MM24_d N_MM24@2_d N_MM25@2_d N_MM25_d N_Q_1
+ N_Q_18 N_Q_17 N_Q_2 N_Q_13 N_Q_16 N_Q_14 N_Q_15 N_Q_19 N_Q_4 N_Q_3
+ PM_DLLx2_ASAP7_75t_R%Q
cc_94 N_Q_1 N_NET085_14 0.000493336f
cc_95 N_Q_18 N_NET085_16 0.000571984f
cc_96 N_Q_17 N_NET085_17 0.000612491f
cc_97 N_Q_2 N_NET085_14 0.00266371f
cc_98 N_Q_13 N_MH_23 0.000301921f
cc_99 N_Q_16 N_MM25@2_g 0.0157914f
cc_100 N_Q_14 N_MM25@2_g 0.0534864f
cc_101 N_Q_15 N_MM25_g 0.0156646f
cc_102 N_Q_19 N_MH_23 0.0068099f
cc_103 N_Q_4 N_MH_2 0.000904046f
cc_104 N_Q_2 N_MM25_g 0.00110289f
cc_105 N_Q_1 N_MM25_g 0.00114323f
cc_106 N_Q_17 N_MH_23 0.0012022f
cc_107 N_Q_4 N_MM25@2_g 0.00122553f
cc_108 N_Q_3 N_MM25@2_g 0.00128925f
cc_109 N_Q_18 N_MH_23 0.00129657f
cc_110 N_Q_18 N_MH_27 0.00215496f
cc_111 N_Q_16 N_MH_2 0.00368597f
cc_112 N_Q_13 N_MM25_g 0.0539698f
x_PM_DLLx2_ASAP7_75t_R%CLKN VSS N_MM22_g N_MM10_g N_MM20_d N_MM21_d N_CLKN_6
+ N_CLKN_5 N_CLKN_23 N_CLKN_13 N_CLKN_14 N_CLKN_1 N_CLKN_16 N_CLKN_18 N_CLKN_19
+ N_CLKN_17 N_CLKN_27 N_CLKN_25 N_CLKN_15 N_CLKN_21 N_CLKN_20 N_CLKN_26
+ N_CLKN_2 PM_DLLx2_ASAP7_75t_R%CLKN
cc_113 N_CLKN_6 N_MM20_g 0.00106627f
cc_114 N_CLKN_5 N_MM20_g 0.00109503f
cc_115 N_CLKN_23 N_MM20_g 0.000248526f
cc_116 N_CLKN_13 N_MM20_g 0.0112204f
cc_117 N_CLKN_14 N_MM20_g 0.0113266f
cc_118 N_CLKN_1 N_CLK_8 0.000419445f
cc_119 N_CLKN_16 N_CLK_8 0.000473525f
cc_120 N_CLKN_18 N_CLK_6 0.000686972f
cc_121 N_CLKN_23 N_CLK_1 0.000776704f
cc_122 N_CLKN_23 N_CLK_4 0.00130371f
cc_123 N_CLKN_19 N_CLK_7 0.0015348f
cc_124 N_CLKN_17 N_CLK_5 0.00177807f
cc_125 N_CLKN_27 N_CLK_8 0.0020032f
cc_126 N_CLKN_25 N_CLK_6 0.0023102f
cc_127 N_CLKN_15 N_CLK_7 0.00242416f
cc_128 N_CLKN_1 N_CLK_1 0.0025247f
cc_129 N_CLKN_19 N_CLK_8 0.00264381f
cc_130 N_CLKN_23 N_CLK_8 0.00323659f
cc_131 N_MM22_g N_MM20_g 0.03533f
x_PM_DLLx2_ASAP7_75t_R%CLKB VSS N_MM1_g N_MM9_g N_MM23_d N_MM22_d N_CLKB_14
+ N_CLKB_5 N_CLKB_17 N_CLKB_4 N_CLKB_16 N_CLKB_21 N_CLKB_6 N_CLKB_15 N_CLKB_19
+ N_CLKB_18 N_CLKB_23 N_CLKB_2 N_CLKB_1 N_CLKB_22 N_CLKB_20
+ PM_DLLx2_ASAP7_75t_R%CLKB
cc_132 N_CLKB_14 N_CLK_5 8.44639e-20
cc_133 N_CLKB_5 N_CLK_5 0.00031786f
cc_134 N_CLKB_17 N_CLK_5 0.000160324f
cc_135 N_CLKB_4 N_CLK_5 0.000435192f
cc_136 N_CLKB_17 N_CLK_6 0.00106721f
cc_137 N_CLKB_16 N_CLK_5 0.00219623f
cc_138 N_CLKB_4 N_MM22_g 0.000858601f
cc_139 N_CLKB_21 N_MM22_g 0.000111867f
cc_140 N_CLKB_6 N_MM10_g 0.000169849f
cc_141 N_CLKB_15 N_MM22_g 0.0111469f
cc_142 N_CLKB_5 N_CLKN_25 0.000336745f
cc_143 N_CLKB_5 N_CLKN_1 0.00039569f
cc_144 N_CLKB_19 N_CLKN_27 0.000404678f
cc_145 N_CLKB_18 N_CLKN_20 0.00151691f
cc_146 N_CLKB_18 N_CLKN_19 0.000473746f
cc_147 N_CLKB_16 N_CLKN_26 0.000582142f
cc_148 N_CLKB_18 N_CLKN_27 0.000628391f
cc_149 N_CLKB_23 N_CLKN_21 0.000645472f
cc_150 N_CLKB_2 N_MM10_g 0.000669269f
cc_151 N_CLKB_1 N_CLKN_2 0.00215049f
cc_152 N_CLKB_15 N_CLKN_1 0.000897935f
cc_153 N_CLKB_5 N_MM22_g 0.00117264f
cc_154 N_MM1_g N_MM10_g 0.00162483f
cc_155 N_CLKB_18 N_CLKN_26 0.00421124f
cc_156 N_CLKB_19 N_CLKN_21 0.00457912f
cc_157 N_CLKB_17 N_CLKN_25 0.00559973f
cc_158 N_MM9_g N_MM10_g 0.00910793f
cc_159 N_CLKB_23 N_CLKN_27 0.0188838f
cc_160 N_CLKB_14 N_MM22_g 0.0389514f
cc_161 N_CLKB_18 N_D_4 0.00352938f
cc_162 N_CLKB_21 N_D_5 0.000890482f
cc_163 N_CLKB_22 N_D_6 0.00089908f
cc_164 N_CLKB_23 N_D_6 0.000906645f
cc_165 N_CLKB_1 N_D_1 0.00273325f
cc_166 N_MM1_g N_MM3_g 0.00506699f
cc_167 N_CLKB_19 N_D_4 0.00921281f
x_PM_DLLx2_ASAP7_75t_R%MH VSS N_MM7_g N_MM25_g N_MM25@2_g N_MM4_d N_MM9_d
+ N_MM1_d N_MM10_d N_MH_22 N_MH_5 N_MH_17 N_MH_19 N_MH_16 N_MH_25 N_MH_27
+ N_MH_20 N_MH_21 N_MH_18 N_MH_6 N_MH_14 N_MH_15 N_MH_26 N_MH_1 N_MH_23 N_MH_2
+ N_MH_24 PM_DLLx2_ASAP7_75t_R%MH
cc_168 N_MH_22 N_MM10_g 0.000139334f
cc_169 N_MH_5 N_CLKN_21 0.000143656f
cc_170 N_MH_17 N_MM10_g 0.000177764f
cc_171 N_MH_19 N_CLKN_21 0.000235268f
cc_172 N_MH_16 N_MM10_g 0.0167259f
cc_173 N_MH_25 N_CLKN_21 0.00053907f
cc_174 N_MH_27 N_CLKN_27 0.000657255f
cc_175 N_MH_5 N_CLKN_2 0.000734988f
cc_176 N_MH_20 N_CLKN_21 0.000815501f
cc_177 N_MH_21 N_CLKN_21 0.00597842f
cc_178 N_MH_18 N_CLKN_27 0.000969597f
cc_179 N_MH_18 N_CLKN_21 0.00103345f
cc_180 N_MH_6 N_MM10_g 0.00110624f
cc_181 N_MH_5 N_MM10_g 0.00138094f
cc_182 N_MH_16 N_CLKN_2 0.00168951f
cc_183 N_MH_14 N_MM10_g 0.0535369f
cc_184 N_MH_14 N_CLKB_20 0.000112131f
cc_185 N_MH_18 N_CLKB_19 0.00134436f
cc_186 N_MH_17 N_MM1_g 0.000151732f
cc_187 N_MH_15 N_MM9_g 0.000170254f
cc_188 N_MH_5 N_CLKB_19 0.00152621f
cc_189 N_MH_20 N_CLKB_20 0.000249869f
cc_190 N_MH_16 N_MM1_g 0.0345563f
cc_191 N_MH_5 N_CLKB_1 0.000269762f
cc_192 N_MH_26 N_CLKB_20 0.000306266f
cc_193 N_MH_1 N_CLKB_6 0.00178859f
cc_194 N_MH_21 N_CLKB_23 0.000620396f
cc_195 N_MH_6 N_MM9_g 0.000632718f
cc_196 N_MH_27 N_CLKB_20 0.00070198f
cc_197 N_MH_22 N_CLKB_6 0.000717063f
cc_198 N_MH_16 N_CLKB_1 0.000794903f
cc_199 N_MH_21 N_CLKB_2 0.000887994f
cc_200 N_MH_5 N_MM1_g 0.00175046f
cc_201 N_MH_21 N_CLKB_20 0.00226127f
cc_202 N_MH_22 N_CLKB_20 0.00405999f
cc_203 N_MH_27 N_CLKB_23 0.00467397f
cc_204 N_MH_18 N_CLKB_23 0.00553462f
cc_205 N_MM7_g N_CLKB_6 0.00635813f
cc_206 N_MH_14 N_MM9_g 0.036925f
cc_207 N_MH_23 N_MM11_g 0.000100265f
cc_208 N_MH_22 N_MM11_g 0.000127807f
cc_209 N_MH_14 N_MM11_g 0.000168215f
cc_210 N_MH_2 N_MM11_g 0.000202436f
cc_211 N_MM7_g N_NET085_10 0.00685f
cc_212 N_MM7_g N_NET085_11 0.00678039f
cc_213 N_MM7_g N_NET085_3 0.000354755f
cc_214 N_MH_27 N_NET085_16 0.000393669f
cc_215 N_MH_6 N_NET085_1 0.000445266f
cc_216 N_MH_22 N_NET085_13 0.000654346f
cc_217 N_MH_1 N_NET085_14 0.000742071f
cc_218 N_MH_22 N_NET085_1 0.000804847f
cc_219 N_MH_1 N_MM11_g 0.000910795f
cc_220 N_MH_24 N_NET085_15 0.000915448f
cc_221 N_MM7_g N_NET085_1 0.001082f
cc_222 N_MH_27 N_NET085_14 0.00268681f
cc_223 N_MH_22 N_NET085_12 0.00304595f
cc_224 N_MH_22 N_NET085_14 0.00367031f
cc_225 N_MH_20 N_NET085_12 0.00367248f
cc_226 N_MM7_g N_MM11_g 0.0288515f
*END of DLLx2_ASAP7_75t_R.pxi
.ENDS
** Design:	DLLx3_ASAP7_75t_R
* Created:	"Fri Aug 17 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "DLLx3_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "DLLx3_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_DLLx3_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00425642f
.ends

.subckt PM_DLLx3_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00432997f
.ends

.subckt PM_DLLx3_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.00552436f
.ends

.subckt PM_DLLx3_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.00550184f
.ends

.subckt PM_DLLx3_ASAP7_75t_R%Q VSS 33 24 25 37 45 48 49 13 3 4 19 18 17 1 2 16
+ 15 14
c1 1 VSS 0.0100448f
c2 2 VSS 0.00994268f
c3 3 VSS 0.00708528f
c4 4 VSS 0.00724593f
c5 13 VSS 0.0046098f
c6 14 VSS 0.00345519f
c7 15 VSS 0.00455141f
c8 16 VSS 0.00344182f
c9 17 VSS 0.0110778f
c10 18 VSS 0.011018f
c11 19 VSS 0.00282517f
c12 20 VSS 0.00194505f
c13 21 VSS 0.00192697f
r1 49 47 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.2025 $X2=0.7705 $Y2=0.2025
r2 2 47 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7560 $Y=0.2025 $X2=0.7705 $Y2=0.2025
r3 15 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7415 $Y=0.2025 $X2=0.7560 $Y2=0.2025
r4 48 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.2025 $X2=0.7415 $Y2=0.2025
r5 16 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.2025 $X2=0.8620 $Y2=0.2025
r6 45 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.2025 $X2=0.8495 $Y2=0.2025
r7 2 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7560 $Y=0.2025
+ $X2=0.7560 $Y2=0.2250
r8 4 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.2025
+ $X2=0.8640 $Y2=0.2250
r9 42 43 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.2250 $X2=0.7695 $Y2=0.2250
r10 40 43 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.2250 $X2=0.7695 $Y2=0.2250
r11 38 39 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.2250 $X2=0.8775 $Y2=0.2250
r12 18 38 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.8235
+ $Y=0.2250 $X2=0.8640 $Y2=0.2250
r13 18 40 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.8235
+ $Y=0.2250 $X2=0.7830 $Y2=0.2250
r14 21 35 5.33101 $w=1.53433e-08 $l=3.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8915 $Y=0.2250 $X2=0.8915 $Y2=0.1915
r15 21 39 1.49343 $w=2.00571e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8915 $Y=0.2250 $X2=0.8775 $Y2=0.2250
r16 14 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.0675 $X2=0.8620 $Y2=0.0675
r17 37 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.0675 $X2=0.8495 $Y2=0.0675
r18 34 35 10.2227 $w=1.4e-08 $l=5.13e-08 $layer=M1 $thickness=3.6e-08 $X=0.8915
+ $Y=0.1402 $X2=0.8915 $Y2=0.1915
r19 33 34 5.43547 $w=1.4e-08 $l=2.72e-08 $layer=M1 $thickness=3.6e-08 $X=0.8915
+ $Y=0.1130 $X2=0.8915 $Y2=0.1402
r20 33 32 2.34373 $w=1.4e-08 $l=1.18e-08 $layer=M1 $thickness=3.6e-08 $X=0.8915
+ $Y=0.1130 $X2=0.8915 $Y2=0.1012
r21 19 20 4.03448 $w=1.56667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8915 $Y=0.0720 $X2=0.8915 $Y2=0.0450
r22 19 32 5.8344 $w=1.4e-08 $l=2.92e-08 $layer=M1 $thickness=3.6e-08 $X=0.8915
+ $Y=0.0720 $X2=0.8915 $Y2=0.1012
r23 3 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.0675
+ $X2=0.8640 $Y2=0.0450
r24 20 31 1.49343 $w=2.00571e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8915 $Y=0.0450 $X2=0.8775 $Y2=0.0450
r25 30 31 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8640
+ $Y=0.0450 $X2=0.8775 $Y2=0.0450
r26 29 30 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.8235
+ $Y=0.0450 $X2=0.8640 $Y2=0.0450
r27 28 29 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.0450 $X2=0.8235 $Y2=0.0450
r28 27 28 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7695
+ $Y=0.0450 $X2=0.7830 $Y2=0.0450
r29 26 27 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.0450 $X2=0.7695 $Y2=0.0450
r30 17 26 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.7445
+ $Y=0.0450 $X2=0.7560 $Y2=0.0450
r31 1 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7560 $Y=0.0675
+ $X2=0.7560 $Y2=0.0450
r32 25 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.0675 $X2=0.7705 $Y2=0.0675
r33 1 23 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7560 $Y=0.0675 $X2=0.7705 $Y2=0.0675
r34 13 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7415 $Y=0.0675 $X2=0.7560 $Y2=0.0675
r35 24 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.0675 $X2=0.7415 $Y2=0.0675
.ends

.subckt PM_DLLx3_ASAP7_75t_R%PU1 VSS 2 4 1
c1 1 VSS 0.000985621f
r1 4 3 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3365 $Y2=0.2025
r2 2 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3195 $Y2=0.2025
r3 1 3 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3195 $Y=0.2025 $X2=0.3365 $Y2=0.2025
.ends

.subckt PM_DLLx3_ASAP7_75t_R%CLK VSS 11 3 8 6 1 7 5 4
c1 1 VSS 0.00254244f
c2 3 VSS 0.0597228f
c3 4 VSS 0.000807828f
c4 5 VSS 0.00434168f
c5 6 VSS 0.00416411f
c6 7 VSS 0.00192763f
c7 8 VSS 0.00179487f
r1 6 17 2.40741 $w=2.45e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.1980 $X2=0.1080 $Y2=0.1710
r2 5 15 4.50612 $w=2.06667e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0630 $X2=0.1080 $Y2=0.0990
r3 16 17 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.1710 $X2=0.1080 $Y2=0.1710
r4 8 13 1.35805 $w=2.83333e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1710 $X2=0.0810 $Y2=0.1485
r5 8 16 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1710 $X2=0.0945 $Y2=0.1710
r6 14 15 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.0990 $X2=0.1080 $Y2=0.0990
r7 7 10 0.483592 $w=3.42308e-08 $l=1.87e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0990 $X2=0.0810 $Y2=0.1177
r8 7 14 0.502848 $w=3.43333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0990 $X2=0.0945 $Y2=0.0990
r9 11 12 0.874462 $w=1.3e-08 $l=3.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1227
r10 11 10 0.291487 $w=1.3e-08 $l=1.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1190 $X2=0.0810 $Y2=0.1177
r11 4 12 2.85657 $w=1.3e-08 $l=1.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1227
r12 4 13 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1485
r13 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r14 1 4 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_DLLx3_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.0418034f
.ends

.subckt PM_DLLx3_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.00472145f
.ends

.subckt PM_DLLx3_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.00473352f
.ends

.subckt PM_DLLx3_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.0419915f
.ends

.subckt PM_DLLx3_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.0418785f
.ends

.subckt PM_DLLx3_ASAP7_75t_R%CLKN VSS 11 12 66 68 6 5 23 14 13 1 16 18 19 17 27
+ 25 15 21 20 26 2
c1 1 VSS 0.0016561f
c2 2 VSS 7.20592e-20
c3 5 VSS 0.00762026f
c4 6 VSS 0.00765707f
c5 11 VSS 0.0598752f
c6 12 VSS 0.00454912f
c7 13 VSS 0.00571706f
c8 14 VSS 0.00560224f
c9 15 VSS 0.00501309f
c10 16 VSS 0.00322905f
c11 17 VSS 0.00475992f
c12 18 VSS 0.00473749f
c13 19 VSS 0.000425828f
c14 20 VSS 0.000393384f
c15 21 VSS 0.000810408f
c16 22 VSS 0.00345478f
c17 23 VSS 0.00145357f
c18 24 VSS 0.00369313f
c19 25 VSS 0.00082045f
c20 26 VSS 0.000405043f
c21 27 VSS 0.0139469f
r1 68 67 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r2 14 67 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r3 66 65 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r4 13 65 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r5 6 63 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0550 $Y2=0.2340
r6 5 60 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0550 $Y2=0.0360
r7 62 63 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.2340 $X2=0.0550 $Y2=0.2340
r8 18 62 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0460 $Y2=0.2340
r9 18 24 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0180 $Y2=0.2340
r10 59 60 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0460
+ $Y=0.0360 $X2=0.0550 $Y2=0.0360
r11 17 59 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0460 $Y2=0.0360
r12 17 22 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0180 $Y2=0.0360
r13 12 57 5.63117 $w=1.26721e-07 $l=2e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4050 $Y2=0.1330
r14 24 56 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.2340 $X2=0.0180 $Y2=0.2070
r15 22 55 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.0360 $X2=0.0180 $Y2=0.0630
r16 2 57 6.49795 $w=1.53e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08 $X=0.4050
+ $Y=0.1440 $X2=0.4050 $Y2=0.1330
r17 16 23 3.9134 $w=1.47857e-08 $l=2.25499e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1755 $X2=0.0165 $Y2=0.1530
r18 16 56 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1755 $X2=0.0180 $Y2=0.2070
r19 54 55 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0990 $X2=0.0180 $Y2=0.0630
r20 15 23 3.9134 $w=1.47857e-08 $l=2.25499e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1305 $X2=0.0165 $Y2=0.1530
r21 15 54 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1305 $X2=0.0180 $Y2=0.0990
r22 52 57 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1440
+ $X2=0.4050 $Y2=0.1330
r23 21 52 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1160 $X2=0.4050 $Y2=0.1440
r24 49 50 1.90199 $w=1.38333e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.0255 $Y=0.1530 $X2=0.0345 $Y2=0.1530
r25 23 49 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0165
+ $Y=0.1530 $X2=0.0255 $Y2=0.1530
r26 25 41 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1980 $X2=0.1890 $Y2=0.1755
r27 47 52 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4050 $Y=0.1530
+ $X2=0.4050 $Y2=0.1440
r28 46 47 21.5701 $w=1.3e-08 $l=9.25e-08 $layer=M2 $thickness=3.6e-08 $X=0.3125
+ $Y=0.1530 $X2=0.4050 $Y2=0.1530
r29 45 46 23.0858 $w=1.3e-08 $l=9.9e-08 $layer=M2 $thickness=3.6e-08 $X=0.2135
+ $Y=0.1530 $X2=0.3125 $Y2=0.1530
r30 44 45 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1530 $X2=0.2135 $Y2=0.1530
r31 43 44 18.1888 $w=1.3e-08 $l=7.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.1110
+ $Y=0.1530 $X2=0.1890 $Y2=0.1530
r32 42 43 18.1888 $w=1.3e-08 $l=7.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.0330
+ $Y=0.1530 $X2=0.1110 $Y2=0.1530
r33 42 50 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.0330 $Y=0.1530
+ $X2=0.0345 $Y2=0.1530
r34 27 42 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.0215
+ $Y=0.1530 $X2=0.0330 $Y2=0.1530
r35 40 41 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1575 $X2=0.1890 $Y2=0.1755
r36 20 26 1.49895 $w=1.95333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1485 $X2=0.1890 $Y2=0.1350
r37 20 40 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1485 $X2=0.1890 $Y2=0.1575
r38 20 44 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.1890 $Y=0.1485
+ $X2=0.1890 $Y2=0.1530
r39 26 39 2.6649 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1705 $Y2=0.1350
r40 38 39 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.1545
+ $Y=0.1350 $X2=0.1705 $Y2=0.1350
r41 37 38 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1455
+ $Y=0.1350 $X2=0.1545 $Y2=0.1350
r42 19 37 1.16595 $w=1.3e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1405
+ $Y=0.1350 $X2=0.1455 $Y2=0.1350
r43 35 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1555 $Y=0.1350
+ $X2=0.1545 $Y2=0.1350
r44 34 35 4.72579 $w=1.53e-08 $l=8e-09 $layer=LIG $thickness=4.8e-08 $X=0.1475
+ $Y=0.1350 $X2=0.1555 $Y2=0.1350
r45 32 34 1.73797 $w=1.72143e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1440 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r46 1 32 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.1340
+ $Y=0.1350 $X2=0.1440 $Y2=0.1350
r47 11 1 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1340 $Y2=0.1350
r48 11 34 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r49 6 14 1e-05
r50 5 13 1e-05
.ends

.subckt PM_DLLx3_ASAP7_75t_R%PD1 VSS 7 10 5 4 1
c1 1 VSS 0.00933465f
c2 4 VSS 0.0031526f
c3 5 VSS 0.00186953f
r1 10 9 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r2 8 9 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r3 5 8 0.123457 $w=8.1e-08 $l=1e-08 $layer=N_src_drn $thickness=1e-09 $X=0.3780
+ $Y=0.0675 $X2=0.3880 $Y2=0.0675
r4 4 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3220 $Y2=0.0675
r5 7 4 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r6 1 5 1e-05
.ends

.subckt PM_DLLx3_ASAP7_75t_R%D VSS 9 3 4 6 5 1
c1 1 VSS 0.0069172f
c2 3 VSS 0.0833645f
c3 4 VSS 0.0057404f
c4 5 VSS 0.00685215f
c5 6 VSS 0.00708882f
r1 6 13 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.2340 $X2=0.2970 $Y2=0.2140
r2 12 13 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1735 $X2=0.2970 $Y2=0.2140
r3 11 12 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1735
r4 10 11 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1215 $X2=0.2970 $Y2=0.1350
r5 9 10 1.16595 $w=1.3e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1165 $X2=0.2970 $Y2=0.1215
r6 9 8 1.28254 $w=1.3e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1165 $X2=0.2970 $Y2=0.1110
r7 4 8 8.27824 $w=1.3e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0755 $X2=0.2970 $Y2=0.1110
r8 4 5 8.03069 $w=1.41392e-08 $l=3.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0755 $X2=0.2970 $Y2=0.0360
r9 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r10 1 11 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_DLLx3_ASAP7_75t_R%PD3 VSS 2 4 1
c1 1 VSS 0.000924064f
r1 4 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0405 $X2=0.4905 $Y2=0.0405
r2 2 1 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0405 $X2=0.4735 $Y2=0.0405
r3 1 3 0.62963 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4735 $Y=0.0405 $X2=0.4905 $Y2=0.0405
.ends

.subckt PM_DLLx3_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.0046208f
.ends

.subckt PM_DLLx3_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.00407065f
.ends

.subckt PM_DLLx3_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.0417957f
.ends

.subckt PM_DLLx3_ASAP7_75t_R%PD2 VSS 7 13 4 1 5
c1 1 VSS 0.00738303f
c2 4 VSS 0.00184671f
c3 5 VSS 0.00234391f
r1 13 12 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r2 5 12 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4880 $Y=0.2295 $X2=0.5005 $Y2=0.2295
r3 10 5 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4725
+ $Y=0.2295 $X2=0.4860 $Y2=0.2295
r4 9 10 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4590
+ $Y=0.2295 $X2=0.4725 $Y2=0.2295
r5 8 9 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4455
+ $Y=0.2295 $X2=0.4590 $Y2=0.2295
r6 1 8 6.3496 $w=2.32e-08 $l=1.35e-08 $layer=LISD $thickness=2.7e-08 $X=0.4320
+ $Y=0.2295 $X2=0.4455 $Y2=0.2295
r7 4 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2295 $X2=0.4300 $Y2=0.2295
r8 7 4 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2295 $X2=0.4175 $Y2=0.2295
.ends

.subckt PM_DLLx3_ASAP7_75t_R%CLKB VSS 12 13 71 73 18 5 17 4 16 21 6 15 19 23 2
+ 1 14 22 20
c1 1 VSS 0.000281628f
c2 2 VSS 9.75104e-20
c3 4 VSS 0.00697118f
c4 5 VSS 0.0073176f
c5 6 VSS 0.0049018f
c6 12 VSS 0.00525393f
c7 13 VSS 0.00505909f
c8 14 VSS 0.00644679f
c9 15 VSS 0.00638327f
c10 16 VSS 0.00981283f
c11 17 VSS 0.00822769f
c12 18 VSS 0.00602886f
c13 19 VSS 0.00114427f
c14 20 VSS 0.00151561f
c15 21 VSS 0.00345064f
c16 22 VSS 0.00293063f
c17 23 VSS 0.0108298f
r1 15 5 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1600 $Y2=0.2160
r2 73 15 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r3 14 4 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1600 $Y2=0.0540
r4 71 14 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r5 5 66 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r6 4 63 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r7 2 54 5.67512 $w=2.4e-08 $l=5e-09 $layer=LISD $thickness=4.02632e-08
+ $X=0.4590 $Y=0.1790 $X2=0.4640 $Y2=0.1790
r8 13 2 2.88446 $w=1.16273e-07 $l=4.4e-08 $layer=LIG $thickness=5.16364e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4590 $Y2=0.1790
r9 66 67 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1845 $Y2=0.2340
r10 17 22 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.2340 $X2=0.2430 $Y2=0.2340
r11 17 67 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.1845 $Y2=0.2340
r12 63 64 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1845 $Y2=0.0360
r13 16 21 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.0360 $X2=0.2430 $Y2=0.0360
r14 16 64 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.1845 $Y2=0.0360
r15 52 54 11.0623 $w=2.14976e-08 $l=2.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4845 $Y=0.1790 $X2=0.4640 $Y2=0.1790
r16 51 52 8.84105 $w=2.02e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4995 $Y=0.1790 $X2=0.4845 $Y2=0.1790
r17 6 49 6.18874 $w=2.02e-08 $l=1.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.5025 $Y=0.1790 $X2=0.5130 $Y2=0.1790
r18 6 51 1.76821 $w=2.02e-08 $l=3e-09 $layer=LISD $thickness=2.7e-08 $X=0.5025
+ $Y=0.1790 $X2=0.4995 $Y2=0.1790
r19 22 46 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2430 $Y2=0.2160
r20 21 43 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0360 $X2=0.2430 $Y2=0.0630
r21 47 49 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5130 $Y=0.1845
+ $X2=0.5130 $Y2=0.1790
r22 20 47 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1680 $X2=0.5130 $Y2=0.1845
r23 45 46 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2025 $X2=0.2430 $Y2=0.2160
r24 44 45 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1935 $X2=0.2430 $Y2=0.2025
r25 42 43 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0990 $X2=0.2430 $Y2=0.0630
r26 41 42 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1215 $X2=0.2430 $Y2=0.0990
r27 40 44 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1845 $X2=0.2430 $Y2=0.1935
r28 18 40 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1530 $X2=0.2430 $Y2=0.1845
r29 18 41 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1530 $X2=0.2430 $Y2=0.1215
r30 38 47 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.5130 $Y=0.1890
+ $X2=0.5130 $Y2=0.1845
r31 37 38 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.4770
+ $Y=0.1890 $X2=0.5130 $Y2=0.1890
r32 36 37 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M2 $thickness=3.6e-08 $X=0.4320
+ $Y=0.1890 $X2=0.4770 $Y2=0.1890
r33 35 36 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M2 $thickness=3.6e-08 $X=0.3870
+ $Y=0.1890 $X2=0.4320 $Y2=0.1890
r34 34 35 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1890 $X2=0.3870 $Y2=0.1890
r35 33 34 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1890 $X2=0.3510 $Y2=0.1890
r36 32 33 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1890 $X2=0.2970 $Y2=0.1890
r37 32 40 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.2430 $Y=0.1890
+ $X2=0.2430 $Y2=0.1845
r38 23 32 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.2315
+ $Y=0.1890 $X2=0.2430 $Y2=0.1890
r39 29 34 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.3510 $Y=0.1890
+ $X2=0.3510 $Y2=0.1890
r40 28 29 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1620 $X2=0.3510 $Y2=0.1890
r41 27 28 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1620
r42 19 27 4.4306 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1160 $X2=0.3510 $Y2=0.1350
r43 12 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r44 1 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
.ends

.subckt PM_DLLx3_ASAP7_75t_R%MH VSS 11 12 13 14 77 81 87 91 23 16 18 20 17 26
+ 28 5 21 22 19 6 15 27 1 24 2 25
c1 1 VSS 0.000512396f
c2 2 VSS 0.0138308f
c3 5 VSS 0.00611566f
c4 6 VSS 0.00510415f
c5 11 VSS 0.0369621f
c6 12 VSS 0.0811128f
c7 13 VSS 0.0805004f
c8 14 VSS 0.0800344f
c9 15 VSS 0.00539117f
c10 16 VSS 0.00152309f
c11 17 VSS 0.0057182f
c12 18 VSS 0.00152006f
c13 19 VSS 0.00948376f
c14 20 VSS 0.00411706f
c15 21 VSS 0.00160822f
c16 22 VSS 0.00066262f
c17 23 VSS 0.000565004f
c18 24 VSS 0.00402843f
c19 25 VSS 0.00329351f
c20 26 VSS 9.7071e-20
c21 27 VSS 0.00287888f
c22 28 VSS 0.0187436f
r1 91 90 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r2 89 90 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3880 $Y=0.2295 $X2=0.3925 $Y2=0.2295
r3 17 89 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3760 $Y=0.2295 $X2=0.3880 $Y2=0.2295
r4 18 17 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2295 $X2=0.3760 $Y2=0.2295
r5 85 86 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r6 87 85 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.1890 $X2=0.3635 $Y2=0.1890
r7 17 86 0.185185 $w=5.4e-08 $l=1e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.1890 $X2=0.3680 $Y2=0.1890
r8 14 71 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=0.8370
+ $Y=0.1350 $X2=0.8370 $Y2=0.1360
r9 12 64 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=0.7290
+ $Y=0.1350 $X2=0.7290 $Y2=0.1360
r10 81 80 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r11 79 80 0.166667 $w=2.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4420 $Y=0.0405 $X2=0.4465 $Y2=0.0405
r12 6 79 0.444445 $w=2.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4300 $Y=0.0405 $X2=0.4420 $Y2=0.0405
r13 16 6 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0405 $X2=0.4300 $Y2=0.0405
r14 15 6 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0810 $X2=0.4300 $Y2=0.0810
r15 77 15 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0810 $X2=0.4175 $Y2=0.0810
r16 73 17 15.0298 $w=2.02e-08 $l=2.55e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.3780 $Y=0.2045 $X2=0.3780 $Y2=0.1790
r17 5 54 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2295
+ $X2=0.3780 $Y2=0.2340
r18 5 73 14.7351 $w=2.02e-08 $l=2.5e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.3780 $Y=0.2295 $X2=0.3780 $Y2=0.2045
r19 69 71 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.8245 $Y=0.1360 $X2=0.8370 $Y2=0.1360
r20 68 69 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.8100 $Y=0.1360 $X2=0.8245 $Y2=0.1360
r21 66 68 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7955 $Y=0.1360 $X2=0.8100 $Y2=0.1360
r22 62 64 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7415 $Y=0.1360 $X2=0.7290 $Y2=0.1360
r23 61 62 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7560 $Y=0.1360 $X2=0.7415 $Y2=0.1360
r24 59 61 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7705 $Y=0.1360 $X2=0.7560 $Y2=0.1360
r25 2 50 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7830 $Y=0.1360
+ $X2=0.7830 $Y2=0.1445
r26 2 59 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7830 $Y=0.1360 $X2=0.7705 $Y2=0.1360
r27 2 66 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7830 $Y=0.1360 $X2=0.7955 $Y2=0.1360
r28 13 2 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=0.7830
+ $Y=0.1350 $X2=0.7830 $Y2=0.1360
r29 6 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0405
+ $X2=0.4320 $Y2=0.0360
r30 54 55 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r31 52 55 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r32 19 27 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4320 $Y=0.2340 $X2=0.4590 $Y2=0.2340
r33 19 52 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4050 $Y2=0.2340
r34 24 50 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1085 $X2=0.7830 $Y2=0.1445
r35 20 25 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4320 $Y=0.0360 $X2=0.4590 $Y2=0.0360
r36 27 45 3.01468 $w=1.741e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4590 $Y2=0.2140
r37 48 50 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.7830 $Y=0.1530
+ $X2=0.7830 $Y2=0.1445
r38 47 48 30.8976 $w=1.3e-08 $l=1.325e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.6505 $Y=0.1530 $X2=0.7830 $Y2=0.1530
r39 46 47 35.678 $w=1.3e-08 $l=1.53e-07 $layer=M2 $thickness=3.6e-08 $X=0.4975
+ $Y=0.1530 $X2=0.6505 $Y2=0.1530
r40 28 46 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M2 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1530 $X2=0.4975 $Y2=0.1530
r41 28 41 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4590 $Y=0.1530
+ $X2=0.4590 $Y2=0.1530
r42 25 40 6.51253 $w=1.552e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4590 $Y2=0.0710
r43 44 45 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2015 $X2=0.4590 $Y2=0.2140
r44 43 44 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1825 $X2=0.4590 $Y2=0.2015
r45 42 43 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1635 $X2=0.4590 $Y2=0.1825
r46 41 42 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1530 $X2=0.4590 $Y2=0.1635
r47 22 41 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1420 $X2=0.4590 $Y2=0.1530
r48 22 26 1.38478 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1420 $X2=0.4590 $Y2=0.1310
r49 39 40 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1015 $X2=0.4590 $Y2=0.0710
r50 21 26 2.78392 $w=1.56471e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1140 $X2=0.4590 $Y2=0.1310
r51 21 39 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1140 $X2=0.4590 $Y2=0.1015
r52 26 38 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1310 $X2=0.4860 $Y2=0.1310
r53 37 38 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1310 $X2=0.4860 $Y2=0.1310
r54 23 35 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.5395
+ $Y=0.1310 $X2=0.5660 $Y2=0.1310
r55 23 37 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.5395
+ $Y=0.1310 $X2=0.5130 $Y2=0.1310
r56 1 32 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.5670
+ $Y=0.1310 $X2=0.5670 $Y2=0.1310
r57 1 35 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1310
+ $X2=0.5660 $Y2=0.1310
r58 11 32 0.314665 $w=2.27e-07 $l=4e-09 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5670 $Y=0.1350 $X2=0.5670 $Y2=0.1310
.ends

.subckt PM_DLLx3_ASAP7_75t_R%NET30 VSS 9 38 43 11 16 1 4 14 3 13 15 10 12
c1 1 VSS 0.00286234f
c2 3 VSS 0.00580945f
c3 4 VSS 0.0066675f
c4 9 VSS 0.03754f
c5 10 VSS 0.00328381f
c6 11 VSS 0.00347158f
c7 12 VSS 0.00128578f
c8 13 VSS 0.00862416f
c9 14 VSS 0.00576832f
c10 15 VSS 0.00340901f
c11 16 VSS 0.00666202f
c12 17 VSS 0.0036886f
r1 11 4 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2295 $X2=0.5920 $Y2=0.2295
r2 43 11 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.2295 $X2=0.5795 $Y2=0.2295
r3 4 40 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2295
+ $X2=0.5940 $Y2=0.2340
r4 40 41 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.2340 $X2=0.6075 $Y2=0.2340
r5 16 36 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.2340 $X2=0.6210 $Y2=0.2205
r6 16 41 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.2340 $X2=0.6075 $Y2=0.2340
r7 10 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.0405 $X2=0.5920 $Y2=0.0405
r8 38 10 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0405 $X2=0.5795 $Y2=0.0405
r9 35 36 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.2095 $X2=0.6210 $Y2=0.2205
r10 34 35 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1850 $X2=0.6210 $Y2=0.2095
r11 33 34 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1660 $X2=0.6210 $Y2=0.1850
r12 32 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1525 $X2=0.6210 $Y2=0.1660
r13 31 32 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1310 $X2=0.6210 $Y2=0.1525
r14 30 31 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1095 $X2=0.6210 $Y2=0.1310
r15 29 30 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0935 $X2=0.6210 $Y2=0.1095
r16 28 29 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0720 $X2=0.6210 $Y2=0.0935
r17 14 27 1.50855 $w=1.55e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0495 $X2=0.6210 $Y2=0.0405
r18 14 28 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0495 $X2=0.6210 $Y2=0.0720
r19 3 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0405
+ $X2=0.5940 $Y2=0.0360
r20 17 26 1.50855 $w=1.55e-08 $l=1.42302e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.0315 $X2=0.6075 $Y2=0.0360
r21 17 27 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0315 $X2=0.6210 $Y2=0.0405
r22 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0360 $X2=0.6075 $Y2=0.0360
r23 24 25 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5825
+ $Y=0.0360 $X2=0.5940 $Y2=0.0360
r24 13 15 7.2121 $w=1.41842e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5510 $Y=0.0360 $X2=0.5130 $Y2=0.0360
r25 13 24 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5510
+ $Y=0.0360 $X2=0.5825 $Y2=0.0360
r26 12 22 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0590 $X2=0.5130 $Y2=0.0820
r27 12 15 3.71425 $w=1.68348e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.0590 $X2=0.5130 $Y2=0.0360
r28 1 19 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.5130
+ $Y=0.0820 $X2=0.5130 $Y2=0.0820
r29 1 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.0820
+ $X2=0.5130 $Y2=0.0820
r30 9 19 0.314665 $w=2.27e-07 $l=5.3e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5130 $Y2=0.0820
.ends


*
.SUBCKT DLLx3_ASAP7_75t_R VSS VDD CLK D Q
*
* VSS VSS
* VDD VDD
* CLK CLK
* D D
* Q Q
*
*

MM20 N_MM20_d N_MM20_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM23 N_MM23_d N_MM22_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM10_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM6 N_MM6_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM24 N_MM24_d N_MM25_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@3 N_MM24@3_d N_MM25@3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@2 N_MM24@2_d N_MM25@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM21 N_MM21_d N_MM20_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM22 N_MM22_d N_MM22_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM25 N_MM25_d N_MM25_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@3 N_MM25@3_d N_MM25@3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@2 N_MM25@2_d N_MM25@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "DLLx3_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "DLLx3_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_DLLx3_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_DLLx3_ASAP7_75t_R%noxref_14
cc_1 N_noxref_14_1 N_MM20_g 0.00368255f
cc_2 N_noxref_14_1 N_CLKN_15 0.000314683f
cc_3 N_noxref_14_1 N_CLKN_5 0.000503361f
cc_4 N_noxref_14_1 N_CLKN_13 0.0278142f
x_PM_DLLx3_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_DLLx3_ASAP7_75t_R%noxref_15
cc_5 N_noxref_15_1 N_MM20_g 0.00367634f
cc_6 N_noxref_15_1 N_CLKN_16 0.000197889f
cc_7 N_noxref_15_1 N_CLKN_6 0.000425988f
cc_8 N_noxref_15_1 N_CLKN_14 0.027902f
cc_9 N_noxref_15_1 N_noxref_14_1 0.00203807f
x_PM_DLLx3_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_DLLx3_ASAP7_75t_R%noxref_24
cc_10 N_noxref_24_1 N_MM25@2_g 0.00150424f
cc_11 N_noxref_24_1 N_Q_14 0.0375658f
x_PM_DLLx3_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_DLLx3_ASAP7_75t_R%noxref_25
cc_12 N_noxref_25_1 N_MM25@2_g 0.00149027f
cc_13 N_noxref_25_1 N_Q_16 0.0376675f
cc_14 N_noxref_25_1 N_noxref_24_1 0.00176809f
x_PM_DLLx3_ASAP7_75t_R%Q VSS Q N_MM24_d N_MM24@3_d N_MM24@2_d N_MM25@2_d
+ N_MM25_d N_MM25@3_d N_Q_13 N_Q_3 N_Q_4 N_Q_19 N_Q_18 N_Q_17 N_Q_1 N_Q_2
+ N_Q_16 N_Q_15 N_Q_14 PM_DLLx3_ASAP7_75t_R%Q
cc_15 N_Q_13 N_MH_24 0.000574105f
cc_16 N_Q_13 N_MM25@2_g 0.000929396f
cc_17 N_Q_13 N_MH_2 0.000529144f
cc_18 N_Q_3 N_MM25@2_g 0.000914765f
cc_19 N_Q_4 N_MM25@2_g 0.000948095f
cc_20 N_Q_19 N_MH_2 0.00112103f
cc_21 N_Q_18 N_MH_24 0.00148115f
cc_22 N_Q_18 N_MH_28 0.00148296f
cc_23 N_Q_17 N_MH_24 0.00152325f
cc_24 N_Q_1 N_MM25_g 0.00204558f
cc_25 N_Q_2 N_MM25_g 0.00216536f
cc_26 N_Q_1 N_MH_24 0.00274498f
cc_27 N_Q_16 N_MM25@2_g 0.0150775f
cc_28 N_Q_15 N_MH_2 0.00679375f
cc_29 N_Q_14 N_MM25@2_g 0.0523241f
cc_30 N_Q_15 N_MM25_g 0.0298833f
cc_31 N_Q_13 N_MM25@3_g 0.0371808f
cc_32 N_Q_13 N_MM25_g 0.0690054f
x_PM_DLLx3_ASAP7_75t_R%PU1 VSS N_MM3_d N_MM1_s N_PU1_1 PM_DLLx3_ASAP7_75t_R%PU1
cc_33 N_PU1_1 N_MM3_g 0.0172488f
cc_34 N_PU1_1 N_MM1_g 0.0169837f
x_PM_DLLx3_ASAP7_75t_R%CLK VSS CLK N_MM20_g N_CLK_8 N_CLK_6 N_CLK_1 N_CLK_7
+ N_CLK_5 N_CLK_4 PM_DLLx3_ASAP7_75t_R%CLK
x_PM_DLLx3_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_DLLx3_ASAP7_75t_R%noxref_18
cc_35 N_noxref_18_1 N_MM3_g 0.00135998f
cc_36 N_noxref_18_1 N_CLKB_18 0.000114861f
cc_37 N_noxref_18_1 N_CLKB_14 0.000714717f
cc_38 N_noxref_18_1 N_noxref_16_1 0.00768305f
cc_39 N_noxref_18_1 N_noxref_17_1 0.000465353f
x_PM_DLLx3_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_DLLx3_ASAP7_75t_R%noxref_17
cc_40 N_noxref_17_1 N_MM22_g 0.00405046f
cc_41 N_noxref_17_1 N_CLKB_5 0.00033745f
cc_42 N_noxref_17_1 N_CLKB_15 0.0270227f
cc_43 N_noxref_17_1 N_noxref_16_1 0.00143201f
x_PM_DLLx3_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_DLLx3_ASAP7_75t_R%noxref_16
cc_44 N_noxref_16_1 N_MM22_g 0.00396869f
cc_45 N_noxref_16_1 N_CLKB_4 0.000355281f
cc_46 N_noxref_16_1 N_CLKB_14 0.0270811f
x_PM_DLLx3_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_DLLx3_ASAP7_75t_R%noxref_23
cc_47 N_noxref_23_1 N_CLKB_6 0.000605151f
cc_48 N_noxref_23_1 N_MM25_g 0.00152968f
cc_49 N_noxref_23_1 N_noxref_20_1 0.000467883f
cc_50 N_noxref_23_1 N_noxref_21_1 0.00759757f
cc_51 N_noxref_23_1 N_noxref_22_1 0.00123263f
x_PM_DLLx3_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_DLLx3_ASAP7_75t_R%noxref_19
cc_52 N_noxref_19_1 N_MM3_g 0.00136904f
cc_53 N_noxref_19_1 N_CLKB_18 0.000108724f
cc_54 N_noxref_19_1 N_CLKB_15 0.000662632f
cc_55 N_noxref_19_1 N_noxref_16_1 0.000464297f
cc_56 N_noxref_19_1 N_noxref_17_1 0.00771177f
cc_57 N_noxref_19_1 N_noxref_18_1 0.00123472f
x_PM_DLLx3_ASAP7_75t_R%CLKN VSS N_MM22_g N_MM10_g N_MM20_d N_MM21_d N_CLKN_6
+ N_CLKN_5 N_CLKN_23 N_CLKN_14 N_CLKN_13 N_CLKN_1 N_CLKN_16 N_CLKN_18 N_CLKN_19
+ N_CLKN_17 N_CLKN_27 N_CLKN_25 N_CLKN_15 N_CLKN_21 N_CLKN_20 N_CLKN_26
+ N_CLKN_2 PM_DLLx3_ASAP7_75t_R%CLKN
cc_58 N_CLKN_6 N_MM20_g 0.00108265f
cc_59 N_CLKN_5 N_MM20_g 0.00110163f
cc_60 N_CLKN_23 N_MM20_g 0.000247314f
cc_61 N_CLKN_14 N_MM20_g 0.0112185f
cc_62 N_CLKN_13 N_MM20_g 0.0112193f
cc_63 N_CLKN_1 N_CLK_8 0.000414216f
cc_64 N_CLKN_16 N_CLK_8 0.000445391f
cc_65 N_CLKN_18 N_CLK_6 0.000742364f
cc_66 N_CLKN_23 N_CLK_1 0.00078207f
cc_67 N_CLKN_19 N_CLK_7 0.00151196f
cc_68 N_CLKN_17 N_CLK_5 0.00184058f
cc_69 N_CLKN_27 N_CLK_8 0.00196324f
cc_70 N_CLKN_23 N_CLK_8 0.00217357f
cc_71 N_CLKN_25 N_CLK_6 0.00233555f
cc_72 N_CLKN_23 N_CLK_4 0.00240868f
cc_73 N_CLKN_15 N_CLK_7 0.0024462f
cc_74 N_CLKN_1 N_CLK_1 0.00254686f
cc_75 N_CLKN_19 N_CLK_8 0.00271284f
cc_76 N_MM22_g N_MM20_g 0.0353094f
x_PM_DLLx3_ASAP7_75t_R%PD1 VSS N_MM5_d N_MM4_s N_PD1_5 N_PD1_4 N_PD1_1
+ PM_DLLx3_ASAP7_75t_R%PD1
cc_77 N_PD1_5 N_CLKN_2 0.000788287f
cc_78 N_PD1_5 N_MM10_g 0.034676f
cc_79 N_PD1_4 N_D_1 0.000679354f
cc_80 N_PD1_4 N_D_4 0.000731415f
cc_81 N_PD1_4 N_MM3_g 0.0358597f
cc_82 N_PD1_4 N_CLKB_19 0.000493819f
cc_83 N_PD1_4 N_CLKB_1 0.00230088f
cc_84 N_PD1_4 N_MM1_g 0.0736833f
cc_85 N_PD1_1 N_MH_20 0.000158206f
cc_86 N_PD1_1 N_MH_6 0.00139015f
cc_87 N_PD1_1 N_MH_15 0.00315833f
x_PM_DLLx3_ASAP7_75t_R%D VSS D N_MM3_g N_D_4 N_D_6 N_D_5 N_D_1
+ PM_DLLx3_ASAP7_75t_R%D
cc_88 N_D_4 N_CLKN_21 0.000139801f
cc_89 N_D_4 N_CLKN_27 0.00281323f
x_PM_DLLx3_ASAP7_75t_R%PD3 VSS N_MM9_s N_MM8_d N_PD3_1 PM_DLLx3_ASAP7_75t_R%PD3
cc_90 N_PD3_1 N_MM9_g 0.0077607f
cc_91 N_PD3_1 N_MM11_g 0.00772875f
x_PM_DLLx3_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_DLLx3_ASAP7_75t_R%noxref_20
cc_92 N_noxref_20_1 N_NET30_10 0.0170504f
cc_93 N_noxref_20_1 N_MM7_g 0.00584493f
x_PM_DLLx3_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_DLLx3_ASAP7_75t_R%noxref_21
cc_94 N_noxref_21_1 N_CLKB_6 0.00286267f
cc_95 N_noxref_21_1 N_NET30_11 0.0163577f
cc_96 N_noxref_21_1 N_MM7_g 0.0052764f
cc_97 N_noxref_21_1 N_noxref_20_1 0.00147867f
x_PM_DLLx3_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_DLLx3_ASAP7_75t_R%noxref_22
cc_98 N_noxref_22_1 N_NET30_10 0.00057376f
cc_99 N_noxref_22_1 N_MM25_g 0.00158224f
cc_100 N_noxref_22_1 N_noxref_20_1 0.00775718f
cc_101 N_noxref_22_1 N_noxref_21_1 0.000450577f
x_PM_DLLx3_ASAP7_75t_R%PD2 VSS N_MM10_s N_MM11_d N_PD2_4 N_PD2_1 N_PD2_5
+ PM_DLLx3_ASAP7_75t_R%PD2
cc_102 N_PD2_4 N_MM10_g 0.0150351f
cc_103 N_PD2_1 N_CLKB_2 0.00101642f
cc_104 N_PD2_5 N_CLKB_6 0.00110067f
cc_105 N_PD2_1 N_MM9_g 0.00216255f
cc_106 N_PD2_5 N_MM9_g 0.00736779f
cc_107 N_PD2_4 N_MM9_g 0.0239933f
cc_108 N_PD2_5 N_MM11_g 0.0147619f
cc_109 N_PD2_1 N_MH_17 0.000614785f
cc_110 N_PD2_1 N_MH_22 0.000390649f
cc_111 N_PD2_1 N_MH_19 0.000404099f
cc_112 N_PD2_4 N_MH_5 0.000590461f
cc_113 N_PD2_1 N_MH_27 0.00210945f
x_PM_DLLx3_ASAP7_75t_R%CLKB VSS N_MM1_g N_MM9_g N_MM23_d N_MM22_d N_CLKB_18
+ N_CLKB_5 N_CLKB_17 N_CLKB_4 N_CLKB_16 N_CLKB_21 N_CLKB_6 N_CLKB_15 N_CLKB_19
+ N_CLKB_23 N_CLKB_2 N_CLKB_1 N_CLKB_14 N_CLKB_22 N_CLKB_20
+ PM_DLLx3_ASAP7_75t_R%CLKB
cc_114 N_CLKB_18 N_CLK_5 0.000107484f
cc_115 N_CLKB_5 N_CLK_5 0.000317164f
cc_116 N_CLKB_17 N_CLK_5 0.000167372f
cc_117 N_CLKB_4 N_CLK_5 0.000440862f
cc_118 N_CLKB_17 N_CLK_6 0.00110334f
cc_119 N_CLKB_16 N_CLK_5 0.00211966f
cc_120 N_CLKB_4 N_MM22_g 0.000876913f
cc_121 N_CLKB_21 N_MM22_g 0.000115182f
cc_122 N_CLKB_6 N_MM10_g 0.00016731f
cc_123 N_CLKB_5 N_CLKN_25 0.000337914f
cc_124 N_CLKB_15 N_MM22_g 0.011286f
cc_125 N_CLKB_5 N_CLKN_1 0.000395894f
cc_126 N_CLKB_19 N_CLKN_27 0.000405046f
cc_127 N_CLKB_18 N_CLKN_20 0.00175835f
cc_128 N_CLKB_18 N_CLKN_19 0.000474463f
cc_129 N_CLKB_16 N_CLKN_26 0.000583127f
cc_130 N_CLKB_18 N_CLKN_27 0.000625888f
cc_131 N_CLKB_23 N_CLKN_21 0.00062891f
cc_132 N_CLKB_2 N_MM10_g 0.000646467f
cc_133 N_CLKB_1 N_CLKN_2 0.00226017f
cc_134 N_CLKB_15 N_CLKN_1 0.000931942f
cc_135 N_CLKB_5 N_MM22_g 0.00122597f
cc_136 N_MM9_g N_MM10_g 0.00368453f
cc_137 N_CLKB_18 N_CLKN_26 0.0041367f
cc_138 N_CLKB_19 N_CLKN_21 0.00462255f
cc_139 N_CLKB_17 N_CLKN_25 0.00571385f
cc_140 N_MM1_g N_MM10_g 0.00705172f
cc_141 N_CLKB_23 N_CLKN_27 0.0187007f
cc_142 N_CLKB_14 N_MM22_g 0.0390121f
cc_143 N_CLKB_19 N_D_4 0.00306465f
cc_144 N_CLKB_22 N_D_6 0.000752931f
cc_145 N_CLKB_23 N_D_6 0.00090171f
cc_146 N_CLKB_21 N_D_5 0.000922394f
cc_147 N_CLKB_1 N_D_1 0.00280096f
cc_148 N_MM1_g N_MM3_g 0.00504648f
cc_149 N_CLKB_18 N_D_4 0.00948655f
x_PM_DLLx3_ASAP7_75t_R%MH VSS N_MM7_g N_MM25_g N_MM25@3_g N_MM25@2_g N_MM4_d
+ N_MM9_d N_MM1_d N_MM10_d N_MH_23 N_MH_16 N_MH_18 N_MH_20 N_MH_17 N_MH_26
+ N_MH_28 N_MH_5 N_MH_21 N_MH_22 N_MH_19 N_MH_6 N_MH_15 N_MH_27 N_MH_1 N_MH_24
+ N_MH_2 N_MH_25 PM_DLLx3_ASAP7_75t_R%MH
cc_150 N_MH_23 N_MM10_g 0.000140642f
cc_151 N_MH_16 N_MM10_g 0.000145946f
cc_152 N_MH_18 N_MM10_g 0.000164091f
cc_153 N_MH_20 N_CLKN_21 0.000225028f
cc_154 N_MH_17 N_MM10_g 0.0166656f
cc_155 N_MH_26 N_CLKN_21 0.000544286f
cc_156 N_MH_28 N_CLKN_27 0.000687636f
cc_157 N_MH_5 N_CLKN_2 0.000776266f
cc_158 N_MH_21 N_CLKN_21 0.000807591f
cc_159 N_MH_22 N_CLKN_21 0.00608403f
cc_160 N_MH_19 N_CLKN_27 0.000958725f
cc_161 N_MH_19 N_CLKN_21 0.00105473f
cc_162 N_MH_6 N_MM10_g 0.00112708f
cc_163 N_MH_5 N_MM10_g 0.00138526f
cc_164 N_MH_17 N_CLKN_2 0.00182607f
cc_165 N_MH_15 N_MM10_g 0.0535464f
cc_166 N_MH_15 N_CLKB_20 0.000110381f
cc_167 N_MH_19 N_CLKB_19 0.00148336f
cc_168 N_MH_18 N_MM1_g 0.000159181f
cc_169 N_MH_16 N_MM9_g 0.000162247f
cc_170 N_MH_5 N_CLKB_19 0.00148505f
cc_171 N_MH_21 N_CLKB_20 0.000265549f
cc_172 N_MH_5 N_CLKB_1 0.000276408f
cc_173 N_MH_17 N_MM1_g 0.0345144f
cc_174 N_MH_27 N_CLKB_20 0.000363683f
cc_175 N_MH_22 N_CLKB_23 0.000453837f
cc_176 N_MH_1 N_CLKB_6 0.00180143f
cc_177 N_MH_6 N_MM9_g 0.0006467f
cc_178 N_MH_28 N_CLKB_20 0.000694889f
cc_179 N_MH_23 N_CLKB_6 0.000716999f
cc_180 N_MH_17 N_CLKB_1 0.000795133f
cc_181 N_MH_22 N_CLKB_2 0.000917262f
cc_182 N_MH_5 N_MM1_g 0.00175828f
cc_183 N_MH_22 N_CLKB_20 0.00214413f
cc_184 N_MH_23 N_CLKB_20 0.00404375f
cc_185 N_MH_28 N_CLKB_23 0.00428303f
cc_186 N_MH_19 N_CLKB_23 0.00550643f
cc_187 N_MM7_g N_CLKB_6 0.00630158f
cc_188 N_MH_15 N_MM9_g 0.0369844f
cc_189 N_MH_20 N_MM11_g 6.26643e-20
cc_190 N_MH_24 N_MM11_g 0.000118984f
cc_191 N_MH_2 N_MM11_g 0.00015832f
cc_192 N_MH_15 N_MM11_g 0.000164913f
cc_193 N_MH_23 N_MM11_g 0.000165815f
cc_194 N_MM7_g N_NET30_11 0.00669456f
cc_195 N_MM7_g N_NET30_3 0.000357037f
cc_196 N_MH_28 N_NET30_16 0.000434769f
cc_197 N_MH_6 N_NET30_1 0.000441714f
cc_198 N_MH_23 N_NET30_13 0.000630777f
cc_199 N_MH_1 N_NET30_14 0.000672862f
cc_200 N_MH_23 N_NET30_1 0.000805663f
cc_201 N_MH_1 N_MM11_g 0.000936853f
cc_202 N_MH_25 N_NET30_15 0.000938748f
cc_203 N_MM7_g N_NET30_1 0.00108204f
cc_204 N_MM7_g N_NET30_10 0.00650399f
cc_205 N_MH_28 N_NET30_14 0.00274986f
cc_206 N_MH_23 N_NET30_12 0.00303406f
cc_207 N_MH_21 N_NET30_12 0.00374374f
cc_208 N_MH_23 N_NET30_14 0.00380377f
cc_209 N_MM7_g N_MM11_g 0.0290045f
x_PM_DLLx3_ASAP7_75t_R%NET30 VSS N_MM11_g N_MM6_d N_MM7_d N_NET30_11 N_NET30_16
+ N_NET30_1 N_NET30_4 N_NET30_14 N_NET30_3 N_NET30_13 N_NET30_15 N_NET30_10
+ N_NET30_12 PM_DLLx3_ASAP7_75t_R%NET30
cc_210 N_MM11_g N_CLKB_2 0.000138371f
cc_211 N_MM11_g N_CLKB_6 0.00514164f
cc_212 N_MM11_g N_CLKB_23 0.000184979f
cc_213 N_MM11_g N_CLKB_20 0.000261132f
cc_214 N_NET30_11 N_CLKB_6 0.000382255f
cc_215 N_NET30_16 N_CLKB_6 0.000391864f
cc_216 N_NET30_1 N_MM9_g 0.000415192f
cc_217 N_NET30_4 N_CLKB_6 0.000848228f
cc_218 N_NET30_14 N_CLKB_6 0.00133086f
cc_219 N_MM11_g N_MM9_g 0.014512f
*END of DLLx3_ASAP7_75t_R.pxi
.ENDS
*
.SUBCKT Comparator A[63] A[62] A[61] A[60] A[59] A[58] A[57] A[56] A[55] A[54] A[53] A[52] A[51] A[50] A[49] A[48] A[47] A[46] A[45] A[44] A[43] A[42] A[41] A[40] A[39] A[38] A[37] A[36] A[35] A[34] A[33] A[32] A[31] A[30] A[29] A[28] A[27] A[26] A[25] A[24] A[23] A[22] A[21] A[20] A[19] A[18] A[17] A[16] A[15] A[14] A[13] A[12] A[11] A[10] A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] B[63] B[62] B[61] B[60] B[59] B[58] B[57] B[56] B[55] B[54] B[53] B[52] B[51] B[50] B[49] B[48] B[47] B[46] B[45] B[44] B[43] B[42] B[41] B[40] B[39] B[38] B[37] B[36] B[35] B[34] B[33] B[32] B[31] B[30] B[29] B[28] B[27] B[26] B[25] B[24] B[23] B[22] B[21] B[20] B[19] B[18] B[17] B[16] B[15] B[14] B[13] B[12] B[11] B[10] B[9] B[8] B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] Out
XU10 n1 n2 n3 n4 n5 Out NOR5xp2_ASAP7_75t_R
XU11 n6 n7 n8 n9 n10 n5 NAND5xp2_ASAP7_75t_R
XU12 B[4] A[4] n14 XOR2xp5_ASAP7_75t_R
XU13 B[5] A[5] n13 XOR2xp5_ASAP7_75t_R
XU14 B[6] A[6] n12 XOR2xp5_ASAP7_75t_R
XU15 B[7] A[7] n11 XOR2xp5_ASAP7_75t_R
XU16 B[3] A[3] n9 XNOR2xp5_ASAP7_75t_R
XU17 B[2] A[2] n8 XNOR2xp5_ASAP7_75t_R
XU18 B[1] A[1] n7 XNOR2xp5_ASAP7_75t_R
XU19 B[0] A[0] n6 XNOR2xp5_ASAP7_75t_R
XU20 n15 n16 n17 n18 n19 n4 NAND5xp2_ASAP7_75t_R
XU21 B[14] A[14] n23 XOR2xp5_ASAP7_75t_R
XU22 B[15] A[15] n22 XOR2xp5_ASAP7_75t_R
XU23 B[8] A[8] n21 XOR2xp5_ASAP7_75t_R
XU24 B[9] A[9] n20 XOR2xp5_ASAP7_75t_R
XU25 B[13] A[13] n18 XNOR2xp5_ASAP7_75t_R
XU26 B[12] A[12] n17 XNOR2xp5_ASAP7_75t_R
XU27 B[11] A[11] n16 XNOR2xp5_ASAP7_75t_R
XU28 B[10] A[10] n15 XNOR2xp5_ASAP7_75t_R
XU29 n24 n25 n26 n27 n28 n3 NAND5xp2_ASAP7_75t_R
XU30 B[20] A[20] n32 XOR2xp5_ASAP7_75t_R
XU31 B[21] A[21] n31 XOR2xp5_ASAP7_75t_R
XU32 B[22] A[22] n30 XOR2xp5_ASAP7_75t_R
XU33 B[23] A[23] n29 XOR2xp5_ASAP7_75t_R
XU34 B[19] A[19] n27 XNOR2xp5_ASAP7_75t_R
XU35 B[18] A[18] n26 XNOR2xp5_ASAP7_75t_R
XU36 B[17] A[17] n25 XNOR2xp5_ASAP7_75t_R
XU37 B[16] A[16] n24 XNOR2xp5_ASAP7_75t_R
XU38 n33 n34 n35 n36 n37 n2 NAND5xp2_ASAP7_75t_R
XU39 B[36] A[36] n41 XOR2xp5_ASAP7_75t_R
XU40 B[37] A[37] n40 XOR2xp5_ASAP7_75t_R
XU41 B[38] A[38] n39 XOR2xp5_ASAP7_75t_R
XU42 B[39] A[39] n38 XOR2xp5_ASAP7_75t_R
XU43 B[35] A[35] n36 XNOR2xp5_ASAP7_75t_R
XU44 B[34] A[34] n35 XNOR2xp5_ASAP7_75t_R
XU45 B[33] A[33] n34 XNOR2xp5_ASAP7_75t_R
XU46 B[32] A[32] n33 XNOR2xp5_ASAP7_75t_R
XU47 n46 n47 n48 n49 n50 n45 NOR5xp2_ASAP7_75t_R
XU48 B[24] A[24] n50 XOR2xp5_ASAP7_75t_R
XU49 B[25] A[25] n49 XOR2xp5_ASAP7_75t_R
XU50 B[26] A[26] n48 XOR2xp5_ASAP7_75t_R
XU51 B[27] A[27] n47 XOR2xp5_ASAP7_75t_R
XU52 B[31] A[31] n54 XNOR2xp5_ASAP7_75t_R
XU53 B[30] A[30] n53 XNOR2xp5_ASAP7_75t_R
XU54 B[29] A[29] n52 XNOR2xp5_ASAP7_75t_R
XU55 B[28] A[28] n51 XNOR2xp5_ASAP7_75t_R
XU56 n55 n56 n57 n58 n59 n44 NOR5xp2_ASAP7_75t_R
XU57 B[56] A[56] n59 XOR2xp5_ASAP7_75t_R
XU58 B[57] A[57] n58 XOR2xp5_ASAP7_75t_R
XU59 B[58] A[58] n57 XOR2xp5_ASAP7_75t_R
XU60 B[59] A[59] n56 XOR2xp5_ASAP7_75t_R
XU61 B[63] A[63] n63 XNOR2xp5_ASAP7_75t_R
XU62 B[62] A[62] n62 XNOR2xp5_ASAP7_75t_R
XU63 B[61] A[61] n61 XNOR2xp5_ASAP7_75t_R
XU64 B[60] A[60] n60 XNOR2xp5_ASAP7_75t_R
XU65 n64 n65 n66 n67 n68 n43 NOR5xp2_ASAP7_75t_R
XU66 B[48] A[48] n68 XOR2xp5_ASAP7_75t_R
XU67 B[49] A[49] n67 XOR2xp5_ASAP7_75t_R
XU68 B[50] A[50] n66 XOR2xp5_ASAP7_75t_R
XU69 B[51] A[51] n65 XOR2xp5_ASAP7_75t_R
XU70 B[55] A[55] n72 XNOR2xp5_ASAP7_75t_R
XU71 B[54] A[54] n71 XNOR2xp5_ASAP7_75t_R
XU72 B[53] A[53] n70 XNOR2xp5_ASAP7_75t_R
XU73 B[52] A[52] n69 XNOR2xp5_ASAP7_75t_R
XU74 n73 n74 n75 n76 n77 n42 NOR5xp2_ASAP7_75t_R
XU75 B[40] A[40] n77 XOR2xp5_ASAP7_75t_R
XU76 B[41] A[41] n76 XOR2xp5_ASAP7_75t_R
XU77 B[42] A[42] n75 XOR2xp5_ASAP7_75t_R
XU78 B[43] A[43] n74 XOR2xp5_ASAP7_75t_R
XU79 B[47] A[47] n81 XNOR2xp5_ASAP7_75t_R
XU80 B[46] A[46] n80 XNOR2xp5_ASAP7_75t_R
XU81 B[45] A[45] n79 XNOR2xp5_ASAP7_75t_R
XU82 B[44] A[44] n78 XNOR2xp5_ASAP7_75t_R
XU83 n42 n43 n44 n45 n1 NAND4xp25_ASAP7_75t_R
XU84 n60 n61 n62 n63 n55 NAND4xp25_ASAP7_75t_R
XU85 n51 n52 n53 n54 n46 NAND4xp25_ASAP7_75t_R
XU86 n69 n70 n71 n72 n64 NAND4xp25_ASAP7_75t_R
XU87 n78 n79 n80 n81 n73 NAND4xp25_ASAP7_75t_R
XU88 n11 n12 n13 n14 n10 NOR4xp25_ASAP7_75t_R
XU89 n20 n21 n22 n23 n19 NOR4xp25_ASAP7_75t_R
XU90 n29 n30 n31 n32 n28 NOR4xp25_ASAP7_75t_R
XU91 n38 n39 n40 n41 n37 NOR4xp25_ASAP7_75t_R
.ENDS



.SUBCKT Adder_4bit A[3] A[2] A[1] A[0] B[3] B[2] B[1] B[0] Output[4] Output[3] Output[2] Output[1] Output[0]
XU3 A[0] B[0] Output[0] XOR2xp5_ASAP7_75t_R
XU4 B[0] A[0] n11 NAND2xp5_ASAP7_75t_R
XU5 B[1] A[1] n11 Output[1] FAx1_ASAP7_75t_R
XU6 B[2] A[2] n6 XNOR2xp5_ASAP7_75t_R
XU7 B[1] A[1] n9 NAND2xp5_ASAP7_75t_R
XU8 n11 n9 n4 NAND2xp5_ASAP7_75t_R
XU9 B[1] A[1] n7 OR2x2_ASAP7_75t_R
XU10 n4 n7 n5 NAND2xp5_ASAP7_75t_R
XU11 n6 n5 Output[2] XOR2xp5_ASAP7_75t_R
XU12 n7 n8 INVx1_ASAP7_75t_R
XU13 B[2] A[2] n10 NAND2xp5_ASAP7_75t_R
XU14 n8 n10 n14 NAND2xp5_ASAP7_75t_R
XU15 B[2] A[2] n13 OR2x2_ASAP7_75t_R
XU16 n11 n10 n9 n12 NAND3xp33_ASAP7_75t_R
XU17 n14 n13 n12 n16 NAND3xp33_ASAP7_75t_R
XU18 B[3] A[3] n15 XNOR2xp5_ASAP7_75t_R
XU19 n16 n15 Output[3] XOR2xp5_ASAP7_75t_R
XU20 n16 n18 INVx1_ASAP7_75t_R
XU21 B[3] A[3] n17 OR2x2_ASAP7_75t_R
XU22 n18 n17 n20 NAND2xp5_ASAP7_75t_R
XU23 B[3] A[3] n19 NAND2xp5_ASAP7_75t_R
XU24 n20 n19 Output[4] NAND2xp5_ASAP7_75t_R
.ENDS



* Design:	AO211x2_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AO211x2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AO211x2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AO211x2_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.00680544f
.ends

.subckt PM_AO211x2_ASAP7_75t_R%NET23 VSS 2 3 1
c1 1 VSS 0.000924087f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_AO211x2_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00563538f
.ends

.subckt PM_AO211x2_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00567272f
.ends

.subckt PM_AO211x2_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.00548431f
.ends

.subckt PM_AO211x2_ASAP7_75t_R%NET20 VSS 19 22 41 42 44 46 1 2 17 13 14 15 3 4
+ 16
c1 1 VSS 0.00793781f
c2 2 VSS 0.00974442f
c3 3 VSS 0.00682849f
c4 4 VSS 0.00555895f
c5 13 VSS 0.00341837f
c6 14 VSS 0.00449947f
c7 15 VSS 0.00323679f
c8 16 VSS 0.00238503f
c9 17 VSS 0.031388f
r1 16 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3760 $Y2=0.2025
r2 46 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r3 44 43 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r4 13 43 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r5 42 40 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r6 2 40 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r7 14 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r8 41 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r9 4 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.2340
r10 1 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0500 $Y2=0.2340
r11 2 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r12 36 37 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3395
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r13 35 36 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2945
+ $Y=0.2340 $X2=0.3395 $Y2=0.2340
r14 34 35 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.2945 $Y2=0.2340
r15 33 34 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r16 29 30 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0590
+ $Y=0.2340 $X2=0.0790 $Y2=0.2340
r17 29 32 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0590
+ $Y=0.2340 $X2=0.0500 $Y2=0.2340
r18 28 30 5.13017 $w=1.3e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1010
+ $Y=0.2340 $X2=0.0790 $Y2=0.2340
r19 27 28 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1255
+ $Y=0.2340 $X2=0.1010 $Y2=0.2340
r20 25 26 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1870 $Y2=0.2340
r21 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r22 24 27 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1255 $Y2=0.2340
r23 23 26 5.13018 $w=1.3e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2090
+ $Y=0.2340 $X2=0.1870 $Y2=0.2340
r24 17 23 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.2335
+ $Y=0.2340 $X2=0.2090 $Y2=0.2340
r25 17 33 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.2335
+ $Y=0.2340 $X2=0.2565 $Y2=0.2340
r26 3 34 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.2340
r27 22 21 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r28 3 21 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r29 18 3 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2600 $Y=0.2025 $X2=0.2720 $Y2=0.2025
r30 15 18 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2600 $Y2=0.2025
r31 19 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r32 1 13 1e-05
.ends

.subckt PM_AO211x2_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.00433792f
.ends

.subckt PM_AO211x2_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.00469537f
.ends

.subckt PM_AO211x2_ASAP7_75t_R%A1 VSS 9 3 4 1 7 6 10
c1 1 VSS 0.00528466f
c2 3 VSS 0.0429698f
c3 4 VSS 0.0432173f
c4 5 VSS 0.00959179f
c5 6 VSS 0.00502857f
c6 7 VSS 0.00232434f
c7 8 VSS 0.0088526f
c8 9 VSS 0.00250953f
c9 10 VSS 0.00434237f
r1 8 27 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0360 $X2=0.0270 $Y2=0.0540
r2 9 6 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1350 $X2=0.0270 $Y2=0.1665
r3 6 10 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1665 $X2=0.0270 $Y2=0.1980
r4 26 27 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0720 $X2=0.0270 $Y2=0.0540
r5 9 5 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1350 $X2=0.0270 $Y2=0.1035
r6 5 26 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1035 $X2=0.0270 $Y2=0.0720
r7 9 24 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1350 $X2=0.0455 $Y2=0.1350
r8 7 22 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.0635
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r9 7 24 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0635
+ $Y=0.1350 $X2=0.0455 $Y2=0.1350
r10 3 17 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0810 $Y2=0.1350
r11 17 18 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0905 $Y2=0.1350
r12 17 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
r13 14 18 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1350 $X2=0.0905 $Y2=0.1350
r14 13 14 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1350 $X2=0.0935 $Y2=0.1350
r15 12 13 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1350 $X2=0.1080 $Y2=0.1350
r16 4 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r17 1 12 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1225 $Y2=0.1350
r18 1 21 3.20232 $w=2.13909e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1460 $Y2=0.1350
r19 4 12 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1225 $Y2=0.1350
r20 4 21 0.905388 $w=2.07755e-07 $l=1.1e-08 $layer=LIG $thickness=5.52727e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1460 $Y2=0.1350
.ends

.subckt PM_AO211x2_ASAP7_75t_R%NET22 VSS 15 18 32 34 13 1 10 11 2 3 12
c1 1 VSS 0.00287279f
c2 2 VSS 0.00390532f
c3 3 VSS 0.00369538f
c4 10 VSS 0.00211008f
c5 11 VSS 0.00216739f
c6 12 VSS 0.00240314f
c7 13 VSS 0.005477f
r1 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2025 $X2=0.5920 $Y2=0.2025
r2 34 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.2025 $X2=0.5795 $Y2=0.2025
r3 32 31 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r4 11 31 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4880 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r5 3 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2025
+ $X2=0.5940 $Y2=0.1980
r6 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2025
+ $X2=0.4900 $Y2=0.1980
r7 28 29 7.22888 $w=1.3e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5630
+ $Y=0.1980 $X2=0.5940 $Y2=0.1980
r8 27 28 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.5335
+ $Y=0.1980 $X2=0.5630 $Y2=0.1980
r9 26 27 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5150
+ $Y=0.1980 $X2=0.5335 $Y2=0.1980
r10 25 26 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.4995
+ $Y=0.1980 $X2=0.5150 $Y2=0.1980
r11 24 25 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4900
+ $Y=0.1980 $X2=0.4995 $Y2=0.1980
r12 23 24 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4810
+ $Y=0.1980 $X2=0.4900 $Y2=0.1980
r13 22 23 10.7267 $w=1.3e-08 $l=4.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.4350
+ $Y=0.1980 $X2=0.4810 $Y2=0.1980
r14 21 22 16.7897 $w=1.3e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.3630
+ $Y=0.1980 $X2=0.4350 $Y2=0.1980
r15 20 21 9.0944 $w=1.3e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1980 $X2=0.3630 $Y2=0.1980
r16 19 20 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3130
+ $Y=0.1980 $X2=0.3240 $Y2=0.1980
r17 13 19 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3105
+ $Y=0.1980 $X2=0.3130 $Y2=0.1980
r18 1 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.1980
r19 18 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r20 16 17 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3340 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r21 1 16 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3220 $Y=0.2025 $X2=0.3340 $Y2=0.2025
r22 10 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3220 $Y2=0.2025
r23 15 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r24 2 11 1e-05
.ends

.subckt PM_AO211x2_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.00536205f
.ends

.subckt PM_AO211x2_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00406618f
.ends

.subckt PM_AO211x2_ASAP7_75t_R%A2 VSS 23 3 4 6 5 10 7 1 8 9
c1 1 VSS 0.0134773f
c2 3 VSS 0.0827318f
c3 4 VSS 0.109538f
c4 5 VSS 0.00171234f
c5 6 VSS 0.00202809f
c6 7 VSS 0.00219522f
c7 8 VSS 0.00198152f
c8 9 VSS 0.00257459f
c9 10 VSS 0.00126829f
r1 6 24 5.75699 $w=1.39091e-08 $l=2.75e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1665 $X2=0.1350 $Y2=0.1390
r2 6 9 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1665 $X2=0.1350 $Y2=0.1980
r3 5 10 5.60393 $w=1.36731e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1035 $X2=0.1350 $Y2=0.1295
r4 5 8 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1035 $X2=0.1350 $Y2=0.0720
r5 23 24 0.561244 $w=1.8e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1335 $X2=0.1350 $Y2=0.1390
r6 23 10 0.408178 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1335 $X2=0.1350 $Y2=0.1295
r7 4 19 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r8 7 21 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r9 23 7 4.24844 $w=9e-09 $l=2.70416e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1335 $X2=0.1620 $Y2=0.1350
r10 17 19 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2305 $Y=0.1350 $X2=0.2430 $Y2=0.1350
r11 16 17 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2160 $Y=0.1350 $X2=0.2305 $Y2=0.1350
r12 15 16 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2015 $Y=0.1350 $X2=0.2160 $Y2=0.1350
r13 13 15 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1985 $Y=0.1350 $X2=0.2015 $Y2=0.1350
r14 12 13 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1985 $Y2=0.1350
r15 12 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
r16 1 12 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1795
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r17 1 14 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.1795
+ $Y=0.1350 $X2=0.1785 $Y2=0.1350
r18 3 12 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1890 $Y2=0.1350
r19 3 14 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.1890 $Y=0.1350 $X2=0.1785 $Y2=0.1350
r20 3 15 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1890 $Y=0.1350 $X2=0.2015 $Y2=0.1350
.ends

.subckt PM_AO211x2_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.0416261f
.ends

.subckt PM_AO211x2_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.0422851f
.ends

.subckt PM_AO211x2_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.0423882f
.ends

.subckt PM_AO211x2_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.0423852f
.ends

.subckt PM_AO211x2_ASAP7_75t_R%Y VSS 21 16 17 28 29 7 10 8 11 1 2
c1 1 VSS 0.0102794f
c2 2 VSS 0.0105868f
c3 7 VSS 0.0045344f
c4 8 VSS 0.00458272f
c5 9 VSS 0.00941892f
c6 10 VSS 0.00960005f
c7 11 VSS 0.00751816f
c8 12 VSS 0.00344242f
c9 13 VSS 0.0034429f
r1 29 27 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.2025 $X2=0.7705 $Y2=0.2025
r2 2 27 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7560 $Y=0.2025 $X2=0.7705 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7415 $Y=0.2025 $X2=0.7560 $Y2=0.2025
r4 28 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.2025 $X2=0.7415 $Y2=0.2025
r5 2 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7560 $Y=0.2025
+ $X2=0.7560 $Y2=0.2340
r6 23 24 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.2340 $X2=0.7965 $Y2=0.2340
r7 10 23 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.7450
+ $Y=0.2340 $X2=0.7560 $Y2=0.2340
r8 13 22 10.0104 $w=1.4764e-08 $l=5e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.2340 $X2=0.8370 $Y2=0.1840
r9 13 24 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8370 $Y=0.2340 $X2=0.7965 $Y2=0.2340
r10 21 22 11.6595 $w=1.3e-08 $l=5e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1340 $X2=0.8370 $Y2=0.1840
r11 11 12 9.77719 $w=1.48e-08 $l=4.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.0850 $X2=0.8370 $Y2=0.0360
r12 21 11 11.4263 $w=1.3e-08 $l=4.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1340 $X2=0.8370 $Y2=0.0850
r13 12 20 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8370 $Y=0.0360 $X2=0.7965 $Y2=0.0360
r14 19 20 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.0360 $X2=0.7965 $Y2=0.0360
r15 18 19 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.7450
+ $Y=0.0360 $X2=0.7560 $Y2=0.0360
r16 9 18 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.7425
+ $Y=0.0360 $X2=0.7450 $Y2=0.0360
r17 1 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7560 $Y=0.0675
+ $X2=0.7560 $Y2=0.0360
r18 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.0675 $X2=0.7705 $Y2=0.0675
r19 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7560 $Y=0.0675 $X2=0.7705 $Y2=0.0675
r20 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7415 $Y=0.0675 $X2=0.7560 $Y2=0.0675
r21 16 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.0675 $X2=0.7415 $Y2=0.0675
.ends

.subckt PM_AO211x2_ASAP7_75t_R%C VSS 5 3 4 7 1 6
c1 1 VSS 0.00788424f
c2 3 VSS 0.0349784f
c3 4 VSS 0.0365674f
c4 5 VSS 0.00398464f
c5 6 VSS 0.00387113f
c6 7 VSS 0.00325083f
r1 7 20 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1620 $X2=0.5130 $Y2=0.1485
r2 6 19 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.0720 $X2=0.5130 $Y2=0.1035
r3 4 16 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1350
r4 5 9 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.1350
+ $X2=0.5130 $Y2=0.1350
r5 5 19 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1035
r6 5 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1485
r7 14 16 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5545 $Y=0.1350 $X2=0.5670 $Y2=0.1350
r8 13 14 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5400 $Y=0.1350 $X2=0.5545 $Y2=0.1350
r9 12 13 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5255 $Y=0.1350 $X2=0.5400 $Y2=0.1350
r10 10 12 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.5225 $Y=0.1350 $X2=0.5255 $Y2=0.1350
r11 9 10 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5225 $Y2=0.1350
r12 1 9 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.5035
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r13 1 11 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.5035
+ $Y=0.1350 $X2=0.5025 $Y2=0.1350
r14 3 9 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r15 3 11 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.5130 $Y=0.1350 $X2=0.5025 $Y2=0.1350
r16 3 12 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5255 $Y2=0.1350
.ends

.subckt PM_AO211x2_ASAP7_75t_R%B VSS 21 3 4 1 5 6 10 8 9
c1 1 VSS 0.00638578f
c2 3 VSS 0.0342605f
c3 4 VSS 0.00805509f
c4 5 VSS 0.00378958f
c5 6 VSS 0.00317452f
c6 7 VSS 0.00327982f
c7 8 VSS 0.00449843f
c8 9 VSS 0.00374239f
c9 10 VSS 0.00256775f
r1 9 25 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1980 $X2=0.2430 $Y2=0.1800
r2 24 25 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1620 $X2=0.2430 $Y2=0.1800
r3 6 10 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.1485 $X2=0.2430 $Y2=0.1350
r4 6 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1485 $X2=0.2430 $Y2=0.1620
r5 5 10 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.1035 $X2=0.2430 $Y2=0.1350
r6 5 8 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.1035 $X2=0.2430 $Y2=0.0720
r7 4 19 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r8 21 7 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2700 $Y2=0.1350
r9 7 10 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2700 $Y=0.1350 $X2=0.2430 $Y2=0.1350
r10 17 19 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3385 $Y=0.1350 $X2=0.3510 $Y2=0.1350
r11 16 17 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3240 $Y=0.1350 $X2=0.3385 $Y2=0.1350
r12 15 16 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3095 $Y=0.1350 $X2=0.3240 $Y2=0.1350
r13 13 15 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.3065 $Y=0.1350 $X2=0.3095 $Y2=0.1350
r14 12 13 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2970
+ $Y=0.1350 $X2=0.3065 $Y2=0.1350
r15 21 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
r16 1 12 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2875
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r17 1 14 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.2875
+ $Y=0.1350 $X2=0.2865 $Y2=0.1350
r18 3 12 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2970 $Y2=0.1350
r19 3 14 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.2970 $Y=0.1350 $X2=0.2865 $Y2=0.1350
r20 3 15 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2970 $Y=0.1350 $X2=0.3095 $Y2=0.1350
.ends

.subckt PM_AO211x2_ASAP7_75t_R%NET014 VSS 15 16 71 73 75 77 80 3 21 17 4 18 24
+ 23 5 19 6 20 27 22 26 28 1 25
c1 1 VSS 0.00853039f
c2 3 VSS 0.00635074f
c3 4 VSS 0.00732125f
c4 5 VSS 0.00706835f
c5 6 VSS 0.00462013f
c6 15 VSS 0.0811757f
c7 16 VSS 0.0808581f
c8 17 VSS 0.00433795f
c9 18 VSS 0.00450228f
c10 19 VSS 0.0044202f
c11 20 VSS 0.00420216f
c12 21 VSS 0.05937f
c13 22 VSS 0.0138926f
c14 23 VSS 0.00394192f
c15 24 VSS 0.00393104f
c16 25 VSS 0.0023374f
c17 26 VSS 0.00289822f
c18 27 VSS 0.000394746f
c19 28 VSS 0.0034956f
r1 80 79 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r2 78 79 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5500 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r3 6 78 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5380 $Y=0.2025 $X2=0.5500 $Y2=0.2025
r4 20 6 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.2025 $X2=0.5380 $Y2=0.2025
r5 77 20 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.2025 $X2=0.5255 $Y2=0.2025
r6 75 74 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r7 17 74 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r8 18 4 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0540 $X2=0.3220 $Y2=0.0540
r9 73 18 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0540 $X2=0.3095 $Y2=0.0540
r10 71 70 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0540 $X2=0.5005 $Y2=0.0540
r11 19 70 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4880 $Y=0.0540 $X2=0.5005 $Y2=0.0540
r12 6 68 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.2025
+ $X2=0.5400 $Y2=0.2340
r13 3 62 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1120 $Y2=0.0360
r14 4 55 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0540
+ $X2=0.3240 $Y2=0.0360
r15 5 52 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0540
+ $X2=0.4900 $Y2=0.0360
r16 68 69 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.2340 $X2=0.5785 $Y2=0.2340
r17 22 28 7.2121 $w=1.41842e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6370 $Y=0.2340 $X2=0.6750 $Y2=0.2340
r18 22 69 13.6416 $w=1.3e-08 $l=5.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.6370
+ $Y=0.2340 $X2=0.5785 $Y2=0.2340
r19 62 63 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1120
+ $Y=0.0360 $X2=0.1305 $Y2=0.0360
r20 61 63 10.0272 $w=1.3e-08 $l=4.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.1735
+ $Y=0.0360 $X2=0.1305 $Y2=0.0360
r21 60 61 8.27824 $w=1.3e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.2090
+ $Y=0.0360 $X2=0.1735 $Y2=0.0360
r22 59 60 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.2335
+ $Y=0.0360 $X2=0.2090 $Y2=0.0360
r23 58 59 11.1931 $w=1.3e-08 $l=4.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2815
+ $Y=0.0360 $X2=0.2335 $Y2=0.0360
r24 56 57 17.7224 $w=1.3e-08 $l=7.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0360 $X2=0.4810 $Y2=0.0360
r25 55 56 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.0360 $X2=0.4050 $Y2=0.0360
r26 54 55 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3130
+ $Y=0.0360 $X2=0.3240 $Y2=0.0360
r27 54 58 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3130
+ $Y=0.0360 $X2=0.2815 $Y2=0.0360
r28 52 53 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4900
+ $Y=0.0360 $X2=0.5085 $Y2=0.0360
r29 52 57 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4900
+ $Y=0.0360 $X2=0.4810 $Y2=0.0360
r30 51 53 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5315
+ $Y=0.0360 $X2=0.5085 $Y2=0.0360
r31 50 51 10.0272 $w=1.3e-08 $l=4.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5745
+ $Y=0.0360 $X2=0.5315 $Y2=0.0360
r32 21 26 7.2121 $w=1.41842e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6370 $Y=0.0360 $X2=0.6750 $Y2=0.0360
r33 21 50 14.5744 $w=1.3e-08 $l=6.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6370
+ $Y=0.0360 $X2=0.5745 $Y2=0.0360
r34 28 49 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.2340 $X2=0.6750 $Y2=0.2160
r35 26 45 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0360 $X2=0.6750 $Y2=0.0540
r36 48 49 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1980 $X2=0.6750 $Y2=0.2160
r37 47 48 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1800 $X2=0.6750 $Y2=0.1980
r38 46 47 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1620 $X2=0.6750 $Y2=0.1800
r39 24 27 2.08435 $w=1.62143e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6750 $Y=0.1480 $X2=0.6750 $Y2=0.1340
r40 24 46 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1480 $X2=0.6750 $Y2=0.1620
r41 44 45 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0720 $X2=0.6750 $Y2=0.0540
r42 23 27 6.04857 $w=1.44516e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6750 $Y=0.1030 $X2=0.6750 $Y2=0.1340
r43 23 44 7.22888 $w=1.3e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1030 $X2=0.6750 $Y2=0.0720
r44 16 37 3.49039 $w=1.235e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=0.7830
+ $Y=0.1350 $X2=0.7830 $Y2=0.1340
r45 25 40 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.1340 $X2=0.7290 $Y2=0.1340
r46 25 27 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7020 $Y=0.1340 $X2=0.6750 $Y2=0.1340
r47 35 37 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7705 $Y=0.1340 $X2=0.7830 $Y2=0.1340
r48 34 35 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7560 $Y=0.1340 $X2=0.7705 $Y2=0.1340
r49 33 34 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7415 $Y=0.1340 $X2=0.7560 $Y2=0.1340
r50 31 33 2.64971 $w=1.44167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.7385 $Y=0.1340 $X2=0.7415 $Y2=0.1340
r51 30 31 3.01694 $w=2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.7290
+ $Y=0.1340 $X2=0.7385 $Y2=0.1340
r52 30 40 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7290 $Y=0.1340
+ $X2=0.7290 $Y2=0.1340
r53 1 30 3.01694 $w=2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.7195
+ $Y=0.1340 $X2=0.7290 $Y2=0.1340
r54 1 32 0.65697 $w=1.665e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.7195
+ $Y=0.1340 $X2=0.7185 $Y2=0.1340
r55 15 30 3.17282 $w=1.28947e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.7290 $Y=0.1350 $X2=0.7290 $Y2=0.1340
r56 15 32 0.812849 $w=2.16824e-07 $l=1.05475e-08 $layer=LIG
+ $thickness=5.5619e-08 $X=0.7290 $Y=0.1350 $X2=0.7185 $Y2=0.1340
r57 15 33 2.80558 $w=1.8426e-07 $l=1.25399e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.7290 $Y=0.1350 $X2=0.7415 $Y2=0.1340
r58 3 17 1e-05
r59 5 19 1e-05
.ends


*
.SUBCKT AO211x2_ASAP7_75t_R VSS VDD A1 A2 B C Y
*
* VSS VSS
* VDD VDD
* A1 A1
* A2 A2
* B B
* C C
* Y Y
*
*

MM24 N_MM24_d N_MM24_g N_MM24_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM5_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM4 N_MM4_d N_MM6_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM8 N_MM8_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8@2 N_MM8@2_d N_MM7@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25 N_MM25_d N_MM25_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@2 N_MM25@2_d N_MM24_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1@2 N_MM1@2_d N_MM1@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@2 N_MM5@2_d N_MM5@2_g N_MM5@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM6_g N_MM6_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6@2 N_MM6@2_d N_MM6@2_g N_MM6@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7@2 N_MM7@2_d N_MM7@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AO211x2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AO211x2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AO211x2_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_AO211x2_ASAP7_75t_R%noxref_19
cc_1 N_noxref_19_1 N_MM6@2_g 0.00155879f
cc_2 N_noxref_19_1 N_NET22_12 0.0360078f
cc_3 N_noxref_19_1 N_noxref_18_1 0.00137616f
x_PM_AO211x2_ASAP7_75t_R%NET23 VSS N_MM24_s N_MM2_d N_NET23_1
+ PM_AO211x2_ASAP7_75t_R%NET23
cc_4 N_NET23_1 N_MM24_g 0.0172721f
cc_5 N_NET23_1 N_MM2_g 0.0173827f
x_PM_AO211x2_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_AO211x2_ASAP7_75t_R%noxref_15
cc_6 N_noxref_15_1 N_MM5@2_g 0.00155091f
cc_7 N_noxref_15_1 N_NET20_16 0.0358597f
cc_8 N_noxref_15_1 N_NET22_10 0.000818016f
cc_9 N_noxref_15_1 N_noxref_14_1 0.00137891f
x_PM_AO211x2_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_AO211x2_ASAP7_75t_R%noxref_13
cc_10 N_noxref_13_1 N_MM25_g 0.00242698f
cc_11 N_noxref_13_1 N_NET20_13 0.0363901f
cc_12 N_noxref_13_1 N_noxref_12_1 0.00191982f
x_PM_AO211x2_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_AO211x2_ASAP7_75t_R%noxref_17
cc_13 N_noxref_17_1 N_MM6_g 0.00156627f
cc_14 N_noxref_17_1 N_NET20_16 0.000544181f
cc_15 N_noxref_17_1 N_NET22_11 0.0362838f
cc_16 N_noxref_17_1 N_noxref_14_1 0.000484578f
cc_17 N_noxref_17_1 N_noxref_15_1 0.00765142f
cc_18 N_noxref_17_1 N_noxref_16_1 0.00136066f
x_PM_AO211x2_ASAP7_75t_R%NET20 VSS N_MM1@2_d N_MM5_s N_MM25@2_d N_MM1_d
+ N_MM25_d N_MM5@2_s N_NET20_1 N_NET20_2 N_NET20_17 N_NET20_13 N_NET20_14
+ N_NET20_15 N_NET20_3 N_NET20_4 N_NET20_16 PM_AO211x2_ASAP7_75t_R%NET20
cc_19 N_NET20_1 N_MM25_g 0.00250531f
cc_20 N_NET20_1 N_A1_6 0.000531487f
cc_21 N_NET20_2 N_MM24_g 0.000748591f
cc_22 N_NET20_17 N_MM24_g 0.00154118f
cc_23 N_NET20_13 N_A1_1 0.00167332f
cc_24 N_NET20_17 N_A1_10 0.00190593f
cc_25 N_NET20_14 N_MM24_g 0.0331569f
cc_26 N_NET20_13 N_MM25_g 0.0355363f
cc_27 N_NET20_15 N_MM2_g 0.000439622f
cc_28 N_NET20_2 N_MM2_g 0.0020884f
cc_29 N_NET20_3 N_MM2_g 0.000730067f
cc_30 N_NET20_15 N_A2_1 0.00145548f
cc_31 N_NET20_17 N_A2_9 0.00485533f
cc_32 N_NET20_15 N_MM1@2_g 0.0331592f
cc_33 N_NET20_14 N_MM2_g 0.0348334f
cc_34 N_NET20_15 N_MM5@2_g 0.000470976f
cc_35 N_NET20_3 N_B_6 0.000592036f
cc_36 N_NET20_4 N_MM5@2_g 0.000946909f
cc_37 N_NET20_3 N_MM5_g 0.00146605f
cc_38 N_NET20_16 N_B_1 0.00164237f
cc_39 N_NET20_17 N_B_9 0.00520133f
cc_40 N_NET20_15 N_MM5_g 0.0332137f
cc_41 N_NET20_16 N_MM5@2_g 0.0352633f
x_PM_AO211x2_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_AO211x2_ASAP7_75t_R%noxref_16
cc_42 N_noxref_16_1 N_MM6_g 0.00354955f
cc_43 N_noxref_16_1 N_NET014_5 0.000381649f
cc_44 N_noxref_16_1 N_NET014_19 0.0270763f
cc_45 N_noxref_16_1 N_NET22_11 0.000586739f
cc_46 N_noxref_16_1 N_noxref_14_1 0.0078905f
cc_47 N_noxref_16_1 N_noxref_15_1 0.000476451f
x_PM_AO211x2_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_AO211x2_ASAP7_75t_R%noxref_12
cc_48 N_noxref_12_1 N_MM25_g 0.0104234f
cc_49 N_noxref_12_1 N_NET014_17 0.000617348f
cc_50 N_noxref_12_1 N_NET20_13 0.000634013f
x_PM_AO211x2_ASAP7_75t_R%A1 VSS A1 N_MM25_g N_MM24_g N_A1_1 N_A1_7 N_A1_6
+ N_A1_10 PM_AO211x2_ASAP7_75t_R%A1
x_PM_AO211x2_ASAP7_75t_R%NET22 VSS N_MM5_d N_MM5@2_d N_MM6_s N_MM6@2_s
+ N_NET22_13 N_NET22_1 N_NET22_10 N_NET22_11 N_NET22_2 N_NET22_3 N_NET22_12
+ PM_AO211x2_ASAP7_75t_R%NET22
cc_51 N_NET22_13 N_MM5@2_g 0.000646821f
cc_52 N_NET22_13 N_B_1 0.00111607f
cc_53 N_NET22_1 N_MM5@2_g 0.00185995f
cc_54 N_NET22_10 N_B_1 0.0024056f
cc_55 N_NET22_10 N_MM5_g 0.0183732f
cc_56 N_NET22_10 N_MM5@2_g 0.0501809f
cc_57 N_NET22_11 N_MM6@2_g 0.000471299f
cc_58 N_NET22_2 N_MM6@2_g 0.00056645f
cc_59 N_NET22_2 N_C 0.000619809f
cc_60 N_NET22_3 N_MM6@2_g 0.00104392f
cc_61 N_NET22_2 N_MM6_g 0.00115303f
cc_62 N_NET22_12 N_C_1 0.00213849f
cc_63 N_NET22_13 N_C_7 0.00555079f
cc_64 N_NET22_11 N_MM6_g 0.0337327f
cc_65 N_NET22_12 N_MM6@2_g 0.0346809f
cc_66 N_NET22_13 N_NET014_20 9.82429e-20
cc_67 N_NET22_13 N_NET014_5 0.000101481f
cc_68 N_NET22_13 N_NET014_23 0.000169836f
cc_69 N_NET22_13 N_NET014_21 0.000170147f
cc_70 N_NET22_13 N_NET014_27 0.000170763f
cc_71 N_NET22_13 N_NET014_6 0.00104209f
cc_72 N_NET22_2 N_NET014_21 0.000406281f
cc_73 N_NET22_13 N_NET014_24 0.000573147f
cc_74 N_NET22_11 N_NET014_20 0.000593702f
cc_75 N_NET22_3 N_NET014_22 0.000616068f
cc_76 N_NET22_12 N_NET014_20 0.00178426f
cc_77 N_NET22_2 N_NET014_6 0.00137186f
cc_78 N_NET22_3 N_NET014_6 0.00514054f
cc_79 N_NET22_13 N_NET014_22 0.0102244f
cc_80 N_NET22_13 N_NET20_4 0.000695583f
cc_81 N_NET22_10 N_NET20_16 0.00181875f
cc_82 N_NET22_1 N_NET20_17 0.000795882f
cc_83 N_NET22_1 N_NET20_3 0.0013626f
cc_84 N_NET22_1 N_NET20_4 0.0052555f
cc_85 N_NET22_13 N_NET20_17 0.010441f
x_PM_AO211x2_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_AO211x2_ASAP7_75t_R%noxref_18
cc_86 N_noxref_18_1 N_MM6@2_g 0.00906645f
cc_87 N_noxref_18_1 N_NET014_21 0.00019555f
cc_88 N_noxref_18_1 N_MM7_g 0.000766948f
cc_89 N_noxref_18_1 N_NET22_12 0.000570202f
x_PM_AO211x2_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_AO211x2_ASAP7_75t_R%noxref_14
cc_90 N_noxref_14_1 N_MM5@2_g 0.00907334f
cc_91 N_noxref_14_1 N_MM6_g 0.000334461f
cc_92 N_noxref_14_1 N_NET014_5 0.000137113f
cc_93 N_noxref_14_1 N_NET014_21 0.000254054f
cc_94 N_noxref_14_1 N_NET014_19 0.00114154f
cc_95 N_noxref_14_1 N_NET20_16 0.000524872f
cc_96 N_noxref_14_1 N_NET22_10 0.000297896f
x_PM_AO211x2_ASAP7_75t_R%A2 VSS A2 N_MM2_g N_MM1@2_g N_A2_6 N_A2_5 N_A2_10
+ N_A2_7 N_A2_1 N_A2_8 N_A2_9 PM_AO211x2_ASAP7_75t_R%A2
cc_97 N_MM2_g N_A1_1 0.000617126f
cc_98 N_MM2_g N_A1_7 0.000620315f
cc_99 N_A2_6 N_A1_7 0.000710933f
cc_100 N_A2_5 N_A1_7 0.000848942f
cc_101 N_A2_10 N_A1_1 0.00156308f
cc_102 N_A2_10 N_A1_7 0.00177906f
cc_103 N_MM2_g N_MM24_g 0.00724199f
x_PM_AO211x2_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_AO211x2_ASAP7_75t_R%noxref_21
cc_104 N_noxref_21_1 N_MM7_g 0.00178463f
cc_105 N_noxref_21_1 N_NET22_12 0.000580327f
cc_106 N_noxref_21_1 N_noxref_18_1 0.000479838f
cc_107 N_noxref_21_1 N_noxref_19_1 0.00765714f
cc_108 N_noxref_21_1 N_noxref_20_1 0.00123817f
x_PM_AO211x2_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_AO211x2_ASAP7_75t_R%noxref_22
cc_109 N_noxref_22_1 N_MM7@2_g 0.00146866f
cc_110 N_noxref_22_1 N_Y_7 0.000840002f
x_PM_AO211x2_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_AO211x2_ASAP7_75t_R%noxref_20
cc_111 N_noxref_20_1 N_MM7_g 0.00186018f
cc_112 N_noxref_20_1 N_noxref_18_1 0.00781908f
x_PM_AO211x2_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_AO211x2_ASAP7_75t_R%noxref_23
cc_113 N_noxref_23_1 N_MM7@2_g 0.00147352f
cc_114 N_noxref_23_1 N_Y_8 0.000846259f
cc_115 N_noxref_23_1 N_noxref_22_1 0.00177282f
x_PM_AO211x2_ASAP7_75t_R%Y VSS Y N_MM8_d N_MM8@2_d N_MM7_d N_MM7@2_d N_Y_7
+ N_Y_10 N_Y_8 N_Y_11 N_Y_1 N_Y_2 PM_AO211x2_ASAP7_75t_R%Y
cc_116 N_Y_7 N_NET014_26 0.000144135f
cc_117 N_Y_7 N_NET014_28 0.000176694f
cc_118 N_Y_7 N_NET014_23 0.00048213f
cc_119 N_Y_7 N_NET014_24 0.000485982f
cc_120 N_Y_7 N_NET014_1 0.00535954f
cc_121 N_Y_10 N_MM7@2_g 0.000609838f
cc_122 N_Y_8 N_MM7@2_g 0.0307345f
cc_123 N_Y_11 N_NET014_1 0.000965903f
cc_124 N_Y_1 N_NET014_25 0.00105263f
cc_125 N_Y_2 N_MM7@2_g 0.0020236f
cc_126 N_Y_1 N_MM7@2_g 0.00212508f
cc_127 N_Y_7 N_MM7_g 0.0372551f
cc_128 N_Y_7 N_MM7@2_g 0.0692846f
x_PM_AO211x2_ASAP7_75t_R%C VSS C N_MM6_g N_MM6@2_g N_C_7 N_C_1 N_C_6
+ PM_AO211x2_ASAP7_75t_R%C
x_PM_AO211x2_ASAP7_75t_R%B VSS B N_MM5_g N_MM5@2_g N_B_1 N_B_5 N_B_6 N_B_10
+ N_B_8 N_B_9 PM_AO211x2_ASAP7_75t_R%B
cc_129 N_B_1 N_MM1@2_g 0.000592689f
cc_130 N_B_5 N_A2_7 0.000662554f
cc_131 N_B_6 N_A2_7 0.000682537f
cc_132 N_B_10 N_A2_1 0.00135524f
cc_133 N_B_10 N_A2_7 0.00191414f
cc_134 N_MM5_g N_MM1@2_g 0.00766064f
x_PM_AO211x2_ASAP7_75t_R%NET014 VSS N_MM7_g N_MM7@2_g N_MM4_d N_MM3_d N_MM24_d
+ N_MM6_d N_MM6@2_d N_NET014_3 N_NET014_21 N_NET014_17 N_NET014_4 N_NET014_18
+ N_NET014_24 N_NET014_23 N_NET014_5 N_NET014_19 N_NET014_6 N_NET014_20
+ N_NET014_27 N_NET014_22 N_NET014_26 N_NET014_28 N_NET014_1 N_NET014_25
+ PM_AO211x2_ASAP7_75t_R%NET014
cc_135 N_NET014_3 N_MM24_g 0.00334752f
cc_136 N_NET014_21 N_MM24_g 0.00144274f
cc_137 N_NET014_17 N_A1_1 0.00247324f
cc_138 N_NET014_17 N_MM25_g 0.0193432f
cc_139 N_NET014_17 N_MM24_g 0.0524644f
cc_140 N_NET014_17 N_A2_8 0.000524861f
cc_141 N_NET014_3 N_A2_8 0.00209999f
cc_142 N_NET014_21 N_A2_7 0.00261071f
cc_143 N_NET014_21 N_A2_8 0.00306344f
cc_144 N_NET014_4 N_MM5@2_g 0.00220531f
cc_145 N_NET014_21 N_MM5@2_g 0.000676564f
cc_146 N_NET014_18 N_B_1 0.000889779f
cc_147 N_NET014_18 N_MM5_g 0.0227428f
cc_148 N_NET014_21 N_B_8 0.0056266f
cc_149 N_NET014_18 N_MM5@2_g 0.029621f
cc_150 N_NET014_24 N_MM6_g 0.0001537f
cc_151 N_NET014_23 N_MM6_g 0.000230717f
cc_152 N_NET014_5 N_MM6_g 0.00142222f
cc_153 N_NET014_19 N_MM6_g 0.0114185f
cc_154 N_NET014_6 N_MM6_g 0.000454361f
cc_155 N_NET014_6 N_C_7 0.00052353f
cc_156 N_NET014_20 N_MM6@2_g 0.0506558f
cc_157 N_NET014_5 N_C 0.000940682f
cc_158 N_NET014_6 N_MM6@2_g 0.00208053f
cc_159 N_NET014_20 N_C_1 0.00283038f
cc_160 N_NET014_21 N_C_6 0.00580566f
cc_161 N_NET014_20 N_MM6_g 0.0330712f
*END of AO211x2_ASAP7_75t_R.pxi
.ENDS
** Design:	AO21x1_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AO21x1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AO21x1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AO21x1_ASAP7_75t_R%NET29 VSS 2 3 1
c1 1 VSS 0.000976561f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_AO21x1_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.00631152f
.ends

.subckt PM_AO21x1_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.0419973f
.ends

.subckt PM_AO21x1_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.00468411f
.ends

.subckt PM_AO21x1_ASAP7_75t_R%A2 VSS 4 3 1
c1 1 VSS 0.00707441f
c2 3 VSS 0.00891636f
c3 4 VSS 0.00524705f
r1 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r2 4 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AO21x1_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00432856f
.ends

.subckt PM_AO21x1_ASAP7_75t_R%B VSS 6 3 4 1
c1 1 VSS 0.00823684f
c2 3 VSS 0.0823832f
c3 4 VSS 0.00441705f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.0980
r2 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AO21x1_ASAP7_75t_R%Y VSS 16 13 22 7 9 2 1 8 10
c1 1 VSS 0.00824904f
c2 2 VSS 0.00744277f
c3 7 VSS 0.0033175f
c4 8 VSS 0.00335708f
c5 9 VSS 0.00586485f
c6 10 VSS 0.00454269f
c7 11 VSS 0.00262028f
r1 9 11 3.36447 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2645 $Y=0.2340 $X2=0.2860 $Y2=0.2340
r2 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2680 $Y2=0.2025
r3 22 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r4 11 20 2.08192 $w=1.85125e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2860 $Y=0.2340 $X2=0.2860 $Y2=0.2180
r5 2 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2765 $Y=0.2025
+ $X2=0.2860 $Y2=0.2000
r6 19 20 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2860
+ $Y=0.2090 $X2=0.2860 $Y2=0.2180
r7 18 19 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2860
+ $Y=0.2000 $X2=0.2860 $Y2=0.2090
r8 17 18 10.7267 $w=1.3e-08 $l=4.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2860
+ $Y=0.1540 $X2=0.2860 $Y2=0.2000
r9 16 17 9.211 $w=1.3e-08 $l=3.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2860
+ $Y=0.1145 $X2=0.2860 $Y2=0.1540
r10 16 15 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2860
+ $Y=0.1145 $X2=0.2860 $Y2=0.0885
r11 14 15 8.04505 $w=1.3e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.2860
+ $Y=0.0540 $X2=0.2860 $Y2=0.0885
r12 10 14 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2860
+ $Y=0.0415 $X2=0.2860 $Y2=0.0540
r13 1 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2765 $Y=0.0675
+ $X2=0.2860 $Y2=0.0540
r14 7 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2680 $Y2=0.0675
r15 13 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
.ends

.subckt PM_AO21x1_ASAP7_75t_R%NET18 VSS 11 20 21 1 7 9 2 8
c1 1 VSS 0.00542855f
c2 2 VSS 0.00728167f
c3 7 VSS 0.00248367f
c4 8 VSS 0.00325045f
c5 9 VSS 0.0121997f
r1 21 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r2 2 19 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r4 20 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r5 2 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r6 15 16 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1235
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r7 14 15 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.0785
+ $Y=0.2340 $X2=0.1235 $Y2=0.2340
r8 13 14 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.0590
+ $Y=0.2340 $X2=0.0785 $Y2=0.2340
r9 12 13 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0500
+ $Y=0.2340 $X2=0.0590 $Y2=0.2340
r10 9 12 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.2340 $X2=0.0500 $Y2=0.2340
r11 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0500 $Y2=0.2340
r12 11 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r13 7 10 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r14 1 7 1e-05
.ends

.subckt PM_AO21x1_ASAP7_75t_R%A1 VSS 10 3 1 6 5 8
c1 1 VSS 0.00248592f
c2 3 VSS 0.0437718f
c3 4 VSS 0.0133284f
c4 5 VSS 0.00399073f
c5 6 VSS 0.00288155f
c6 7 VSS 0.00197868f
c7 8 VSS 0.0033909f
r1 8 16 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1980 $X2=0.0270 $Y2=0.1765
r2 5 7 3.2503 $w=1.53684e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1540 $X2=0.0270 $Y2=0.1350
r3 5 16 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1540 $X2=0.0270 $Y2=0.1765
r4 4 7 7.44771 $w=1.42162e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0980 $X2=0.0270 $Y2=0.1350
r5 7 12 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1350 $X2=0.0455 $Y2=0.1350
r6 10 6 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0635 $Y2=0.1350
r7 6 12 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0635
+ $Y=0.1350 $X2=0.0455 $Y2=0.1350
r8 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r9 10 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AO21x1_ASAP7_75t_R%NET16 VSS 9 39 40 43 44 11 3 12 13 10 4 14 15 1 16
c1 1 VSS 0.00338345f
c2 3 VSS 0.00292f
c3 4 VSS 0.00863649f
c4 9 VSS 0.0797218f
c5 10 VSS 0.00390866f
c6 11 VSS 0.0023921f
c7 12 VSS 0.00289613f
c8 13 VSS 0.00878938f
c9 14 VSS 0.00277014f
c10 15 VSS 0.00285331f
c11 16 VSS 0.000454579f
r1 44 42 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r2 3 42 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r3 11 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r4 43 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
r5 40 38 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r6 4 38 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r7 10 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r8 39 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1475 $Y2=0.0675
r9 3 34 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.1980
r10 4 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0675
+ $X2=0.1620 $Y2=0.0360
r11 34 35 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.1980 $X2=0.1215 $Y2=0.1980
r12 32 35 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1980 $X2=0.1215 $Y2=0.1980
r13 31 32 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1460
+ $Y=0.1980 $X2=0.1350 $Y2=0.1980
r14 30 31 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.1980 $X2=0.1460 $Y2=0.1980
r15 29 30 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.1780
+ $Y=0.1980 $X2=0.1620 $Y2=0.1980
r16 28 29 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1980 $X2=0.1780 $Y2=0.1980
r17 27 28 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2140
+ $Y=0.1980 $X2=0.1890 $Y2=0.1980
r18 12 16 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2320 $Y=0.1980 $X2=0.2430 $Y2=0.1980
r19 12 27 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2320
+ $Y=0.1980 $X2=0.2140 $Y2=0.1980
r20 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r21 23 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r22 13 15 4.55457 $w=1.3814e-08 $l=2.75545e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.0360 $X2=0.2430 $Y2=0.0415
r23 13 23 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r24 16 21 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.1980 $X2=0.2430 $Y2=0.1765
r25 15 20 3.27203 $w=1.40938e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0415 $X2=0.2430 $Y2=0.0575
r26 19 21 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1540 $X2=0.2430 $Y2=0.1765
r27 18 19 4.4306 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1540
r28 14 18 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0980 $X2=0.2430 $Y2=0.1350
r29 14 20 9.44418 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0980 $X2=0.2430 $Y2=0.0575
r30 9 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r31 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends


*
.SUBCKT AO21x1_ASAP7_75t_R VSS VDD A1 A2 B Y
*
* VSS VSS
* VDD VDD
* A1 A1
* A2 A2
* B B
* Y Y
*
*

MM2 N_MM2_d N_MM2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g N_MM3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM2_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM3_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 VDD N_MM4_g N_MM0_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AO21x1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AO21x1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AO21x1_ASAP7_75t_R%NET29 VSS N_MM2_d N_MM3_s N_NET29_1
+ PM_AO21x1_ASAP7_75t_R%NET29
cc_1 N_NET29_1 N_MM2_g 0.0172449f
cc_2 N_NET29_1 N_MM3_g 0.0173677f
x_PM_AO21x1_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_AO21x1_ASAP7_75t_R%noxref_11
cc_3 N_noxref_11_1 N_MM2_g 0.00213692f
cc_4 N_noxref_11_1 N_NET18_7 0.0361475f
cc_5 N_noxref_11_1 N_noxref_10_1 0.00177059f
x_PM_AO21x1_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_AO21x1_ASAP7_75t_R%noxref_10
cc_6 N_noxref_10_1 N_MM2_g 0.00220841f
cc_7 N_noxref_10_1 N_NET18_7 0.000478464f
x_PM_AO21x1_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_AO21x1_ASAP7_75t_R%noxref_12
cc_8 N_noxref_12_1 N_MM7_g 0.00141587f
cc_9 N_noxref_12_1 N_Y_7 0.0390959f
x_PM_AO21x1_ASAP7_75t_R%A2 VSS A2 N_MM3_g N_A2_1 PM_AO21x1_ASAP7_75t_R%A2
cc_10 N_A2_1 N_A1_1 0.00121958f
cc_11 N_A2 N_A1_6 0.00262189f
cc_12 N_MM3_g N_MM2_g 0.00636344f
x_PM_AO21x1_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_AO21x1_ASAP7_75t_R%noxref_13
cc_13 N_noxref_13_1 N_MM7_g 0.00140437f
cc_14 N_noxref_13_1 N_Y_8 0.0393579f
cc_15 N_noxref_13_1 N_noxref_12_1 0.00172546f
x_PM_AO21x1_ASAP7_75t_R%B VSS B N_MM4_g N_B_4 N_B_1 PM_AO21x1_ASAP7_75t_R%B
cc_16 N_B_4 N_A2 0.00328746f
cc_17 N_MM4_g N_MM3_g 0.00491197f
x_PM_AO21x1_ASAP7_75t_R%Y VSS Y N_MM7_d N_MM8_d N_Y_7 N_Y_9 N_Y_2 N_Y_1 N_Y_8
+ N_Y_10 PM_AO21x1_ASAP7_75t_R%Y
cc_18 N_Y_7 N_NET16_15 0.000592823f
cc_19 N_Y_7 N_NET16_1 0.000823471f
cc_20 N_Y_9 N_NET16_12 0.00085593f
cc_21 N_Y_2 N_MM7_g 0.00138923f
cc_22 N_Y_1 N_MM7_g 0.00158938f
cc_23 N_Y_8 N_NET16_1 0.00163043f
cc_24 N_Y_9 N_NET16_16 0.00280552f
cc_25 N_Y_8 N_MM7_g 0.0154172f
cc_26 N_Y_10 N_NET16_14 0.00959809f
cc_27 N_Y_7 N_MM7_g 0.0549478f
x_PM_AO21x1_ASAP7_75t_R%NET18 VSS N_MM1_d N_MM5_d N_MM0_s N_NET18_1 N_NET18_7
+ N_NET18_9 N_NET18_2 N_NET18_8 PM_AO21x1_ASAP7_75t_R%NET18
cc_28 N_NET18_1 N_A1_5 0.000536468f
cc_29 N_NET18_7 N_A1_1 0.000796372f
cc_30 N_NET18_1 N_MM2_g 0.00195287f
cc_31 N_NET18_9 N_A1_8 0.00342356f
cc_32 N_NET18_7 N_MM2_g 0.0350057f
cc_33 N_NET18_2 N_MM3_g 0.00088255f
cc_34 N_NET18_8 N_MM3_g 0.034714f
cc_35 N_NET18_2 N_MM4_g 0.000883302f
cc_36 N_NET18_8 N_MM4_g 0.0347696f
cc_37 N_NET18_7 N_NET16_12 0.000564535f
cc_38 N_NET18_8 N_NET16_11 0.00174589f
cc_39 N_NET18_9 N_NET16_3 0.000765497f
cc_40 N_NET18_1 N_NET16_3 0.00136645f
cc_41 N_NET18_2 N_NET16_3 0.00475932f
cc_42 N_NET18_9 N_NET16_12 0.00980475f
x_PM_AO21x1_ASAP7_75t_R%A1 VSS A1 N_MM2_g N_A1_1 N_A1_6 N_A1_5 N_A1_8
+ PM_AO21x1_ASAP7_75t_R%A1
x_PM_AO21x1_ASAP7_75t_R%NET16 VSS N_MM7_g N_MM3_d N_MM4_d N_MM1_s N_MM5_s
+ N_NET16_11 N_NET16_3 N_NET16_12 N_NET16_13 N_NET16_10 N_NET16_4 N_NET16_14
+ N_NET16_15 N_NET16_1 N_NET16_16 PM_AO21x1_ASAP7_75t_R%NET16
cc_43 N_NET16_11 N_A1_1 0.00123364f
cc_44 N_NET16_3 N_MM2_g 0.000956747f
cc_45 N_NET16_12 N_A1_6 0.00123989f
cc_46 N_NET16_11 N_MM2_g 0.0361568f
cc_47 N_NET16_13 N_A2 0.000534141f
cc_48 N_NET16_3 N_A2_1 0.00059141f
cc_49 N_NET16_3 N_MM3_g 0.000916397f
cc_50 N_NET16_12 N_A2 0.00123608f
cc_51 N_NET16_10 N_A2_1 0.00144569f
cc_52 N_NET16_4 N_MM3_g 0.00159258f
cc_53 N_NET16_4 N_A2 0.00267555f
cc_54 N_NET16_11 N_MM3_g 0.0152218f
cc_55 N_NET16_10 N_MM3_g 0.054948f
cc_56 N_NET16_4 N_MM4_g 0.00195535f
cc_57 N_NET16_13 N_B_4 0.00101398f
cc_58 N_NET16_12 N_B_4 0.0012289f
cc_59 N_NET16_10 N_B_1 0.00125474f
cc_60 N_MM7_g N_MM4_g 0.00162583f
cc_61 N_NET16_14 N_B_4 0.00617909f
cc_62 N_NET16_10 N_MM4_g 0.0372858f
*END of AO21x1_ASAP7_75t_R.pxi
.ENDS
** Design:	AO21x2_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AO21x2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AO21x2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AO21x2_ASAP7_75t_R%NET29 VSS 2 3 1
c1 1 VSS 0.00100533f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_AO21x2_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.00639359f
.ends

.subckt PM_AO21x2_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.0419959f
.ends

.subckt PM_AO21x2_ASAP7_75t_R%A2 VSS 4 3 1
c1 1 VSS 0.00672345f
c2 3 VSS 0.00874682f
c3 4 VSS 0.00499594f
r1 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r2 4 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AO21x2_ASAP7_75t_R%NET18 VSS 11 20 21 1 7 9 2 8
c1 1 VSS 0.00542223f
c2 2 VSS 0.00727752f
c3 7 VSS 0.00248076f
c4 8 VSS 0.00323863f
c5 9 VSS 0.0112495f
r1 21 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r2 2 19 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r4 20 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r5 2 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r6 15 16 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1235
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r7 14 15 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.0785
+ $Y=0.2340 $X2=0.1235 $Y2=0.2340
r8 13 14 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.0590
+ $Y=0.2340 $X2=0.0785 $Y2=0.2340
r9 12 13 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0500
+ $Y=0.2340 $X2=0.0590 $Y2=0.2340
r10 9 12 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.2340 $X2=0.0500 $Y2=0.2340
r11 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0500 $Y2=0.2340
r12 11 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r13 7 10 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r14 1 7 1e-05
.ends

.subckt PM_AO21x2_ASAP7_75t_R%B VSS 6 3 4 1
c1 1 VSS 0.00815315f
c2 3 VSS 0.0823922f
c3 4 VSS 0.00437323f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.0980
r2 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AO21x2_ASAP7_75t_R%A1 VSS 10 3 1 6 5 8
c1 1 VSS 0.00255517f
c2 3 VSS 0.0437697f
c3 4 VSS 0.0134189f
c4 5 VSS 0.00398457f
c5 6 VSS 0.00292619f
c6 7 VSS 0.00201798f
c7 8 VSS 0.0034281f
r1 8 16 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1980 $X2=0.0270 $Y2=0.1765
r2 5 7 3.2503 $w=1.53684e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1540 $X2=0.0270 $Y2=0.1350
r3 5 16 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1540 $X2=0.0270 $Y2=0.1765
r4 4 7 7.44771 $w=1.42162e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0980 $X2=0.0270 $Y2=0.1350
r5 7 12 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1350 $X2=0.0455 $Y2=0.1350
r6 10 6 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0635 $Y2=0.1350
r7 6 12 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0635
+ $Y=0.1350 $X2=0.0455 $Y2=0.1350
r8 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r9 10 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AO21x2_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.0426243f
.ends

.subckt PM_AO21x2_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.0425295f
.ends

.subckt PM_AO21x2_ASAP7_75t_R%Y VSS 22 17 18 32 33 7 9 11 2 1 12 8
c1 1 VSS 0.0130984f
c2 2 VSS 0.00961412f
c3 7 VSS 0.00367395f
c4 8 VSS 0.00445875f
c5 9 VSS 0.00872692f
c6 10 VSS 0.000698455f
c7 11 VSS 0.00583156f
c8 12 VSS 0.00266066f
c9 13 VSS 0.00157276f
c10 14 VSS 0.00317354f
r1 33 31 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r2 2 31 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r4 32 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r5 2 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2685 $Y2=0.2340
r6 25 26 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2775
+ $Y=0.2340 $X2=0.2865 $Y2=0.2340
r7 25 28 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2775
+ $Y=0.2340 $X2=0.2685 $Y2=0.2340
r8 9 14 2.89809 $w=1.53077e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3045 $Y=0.2340 $X2=0.3240 $Y2=0.2340
r9 9 26 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3045
+ $Y=0.2340 $X2=0.2865 $Y2=0.2340
r10 14 24 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.2340 $X2=0.3240 $Y2=0.2160
r11 23 24 12.8254 $w=1.3e-08 $l=5.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1610 $X2=0.3240 $Y2=0.2160
r12 22 23 10.8433 $w=1.3e-08 $l=4.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1145 $X2=0.3240 $Y2=0.1610
r13 22 11 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1145 $X2=0.3240 $Y2=0.1005
r14 11 13 3.59766 $w=1.692e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3240 $Y=0.1005 $X2=0.3240 $Y2=0.0780
r15 10 21 3.36689 $w=1.53077e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3045 $Y=0.0780 $X2=0.2850 $Y2=0.0780
r16 10 13 2.89809 $w=1.53077e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3045 $Y=0.0780 $X2=0.3240 $Y2=0.0780
r17 20 21 1.61797 $w=1.675e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2850 $Y=0.0660 $X2=0.2850 $Y2=0.0780
r18 19 20 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2850
+ $Y=0.0540 $X2=0.2850 $Y2=0.0660
r19 12 19 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2850
+ $Y=0.0415 $X2=0.2850 $Y2=0.0540
r20 1 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2760 $Y=0.0675
+ $X2=0.2850 $Y2=0.0540
r21 18 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r22 1 16 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r23 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r24 17 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
.ends

.subckt PM_AO21x2_ASAP7_75t_R%NET16 VSS 9 10 51 52 55 56 3 12 13 14 4 11 15 16
+ 1 17
c1 1 VSS 0.00780803f
c2 3 VSS 0.00287362f
c3 4 VSS 0.008619f
c4 9 VSS 0.0807431f
c5 10 VSS 0.0807014f
c6 11 VSS 0.00756731f
c7 12 VSS 0.00590907f
c8 13 VSS 0.00453916f
c9 14 VSS 0.0106999f
c10 15 VSS 0.00483495f
c11 16 VSS 0.00268689f
c12 17 VSS 0.000547718f
r1 56 54 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r2 3 54 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r3 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r4 55 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
r5 52 50 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r6 4 50 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r7 11 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r8 51 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1475 $Y2=0.0675
r9 3 46 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.1980
r10 4 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0675
+ $X2=0.1620 $Y2=0.0360
r11 46 47 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.1980 $X2=0.1215 $Y2=0.1980
r12 44 47 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1980 $X2=0.1215 $Y2=0.1980
r13 43 44 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1460
+ $Y=0.1980 $X2=0.1350 $Y2=0.1980
r14 42 43 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.1980 $X2=0.1460 $Y2=0.1980
r15 41 42 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.1780
+ $Y=0.1980 $X2=0.1620 $Y2=0.1980
r16 40 41 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1980 $X2=0.1780 $Y2=0.1980
r17 39 40 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2140
+ $Y=0.1980 $X2=0.1890 $Y2=0.1980
r18 13 17 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2320 $Y=0.1980 $X2=0.2430 $Y2=0.1980
r19 13 39 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2320
+ $Y=0.1980 $X2=0.2140 $Y2=0.1980
r20 37 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r21 35 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r22 14 16 4.55457 $w=1.3814e-08 $l=2.75545e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.0360 $X2=0.2430 $Y2=0.0415
r23 14 35 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r24 17 32 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.1980 $X2=0.2430 $Y2=0.1765
r25 16 31 3.27203 $w=1.40938e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0415 $X2=0.2430 $Y2=0.0575
r26 10 26 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r27 30 31 4.89699 $w=1.3e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0785 $X2=0.2430 $Y2=0.0575
r28 29 32 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1540 $X2=0.2430 $Y2=0.1765
r29 28 29 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1540
r30 15 28 6.64591 $w=1.3e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1065 $X2=0.2430 $Y2=0.1350
r31 15 30 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1065 $X2=0.2430 $Y2=0.0785
r32 24 26 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2845 $Y=0.1350 $X2=0.2970 $Y2=0.1350
r33 23 24 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2700 $Y=0.1350 $X2=0.2845 $Y2=0.1350
r34 22 23 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2555 $Y=0.1350 $X2=0.2700 $Y2=0.1350
r35 20 22 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.2525 $Y=0.1350 $X2=0.2555 $Y2=0.1350
r36 19 20 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2525 $Y2=0.1350
r37 19 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
r38 1 19 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2335
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r39 1 21 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.2335
+ $Y=0.1350 $X2=0.2325 $Y2=0.1350
r40 9 19 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2430 $Y2=0.1350
r41 9 21 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.2430 $Y=0.1350 $X2=0.2325 $Y2=0.1350
r42 9 22 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2555 $Y2=0.1350
.ends


*
.SUBCKT AO21x2_ASAP7_75t_R VSS VDD A1 A2 B Y
*
* VSS VSS
* VDD VDD
* A1 A1
* A2 A2
* B B
* Y Y
*
*

MM2 N_MM2_d N_MM2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g N_MM3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7@2 N_MM7@2_d N_MM7@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM2_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM3_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 VDD N_MM4_g N_MM0_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8@2 N_MM8@2_d N_MM7@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AO21x2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AO21x2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AO21x2_ASAP7_75t_R%NET29 VSS N_MM2_d N_MM3_s N_NET29_1
+ PM_AO21x2_ASAP7_75t_R%NET29
cc_1 N_NET29_1 N_MM2_g 0.0172535f
cc_2 N_NET29_1 N_MM3_g 0.0173304f
x_PM_AO21x2_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_AO21x2_ASAP7_75t_R%noxref_11
cc_3 N_noxref_11_1 N_MM2_g 0.00214264f
cc_4 N_noxref_11_1 N_NET18_7 0.0361174f
cc_5 N_noxref_11_1 N_noxref_10_1 0.00176148f
x_PM_AO21x2_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_AO21x2_ASAP7_75t_R%noxref_10
cc_6 N_noxref_10_1 N_MM2_g 0.00221081f
cc_7 N_noxref_10_1 N_NET18_7 0.000477749f
x_PM_AO21x2_ASAP7_75t_R%A2 VSS A2 N_MM3_g N_A2_1 PM_AO21x2_ASAP7_75t_R%A2
cc_8 N_A2_1 N_A1_1 0.00124777f
cc_9 N_A2 N_A1_6 0.00247978f
cc_10 N_MM3_g N_MM2_g 0.00635824f
x_PM_AO21x2_ASAP7_75t_R%NET18 VSS N_MM1_d N_MM5_d N_MM0_s N_NET18_1 N_NET18_7
+ N_NET18_9 N_NET18_2 N_NET18_8 PM_AO21x2_ASAP7_75t_R%NET18
cc_11 N_NET18_1 N_A1_5 0.000519571f
cc_12 N_NET18_7 N_A1_1 0.00085106f
cc_13 N_NET18_1 N_MM2_g 0.00195059f
cc_14 N_NET18_9 N_A1_8 0.00336041f
cc_15 N_NET18_7 N_MM2_g 0.0349689f
cc_16 N_NET18_2 N_MM3_g 0.00089694f
cc_17 N_NET18_8 N_MM3_g 0.0346579f
cc_18 N_NET18_2 N_MM4_g 0.000904021f
cc_19 N_NET18_8 N_MM4_g 0.034733f
cc_20 N_NET18_7 N_NET16_12 0.000563871f
cc_21 N_NET18_8 N_NET16_12 0.00174161f
cc_22 N_NET18_9 N_NET16_3 0.000764597f
cc_23 N_NET18_1 N_NET16_3 0.00136522f
cc_24 N_NET18_2 N_NET16_3 0.00477953f
cc_25 N_NET18_9 N_NET16_13 0.0100619f
x_PM_AO21x2_ASAP7_75t_R%B VSS B N_MM4_g N_B_4 N_B_1 PM_AO21x2_ASAP7_75t_R%B
cc_26 N_B_4 N_A2 0.0032541f
cc_27 N_MM4_g N_MM3_g 0.00490948f
x_PM_AO21x2_ASAP7_75t_R%A1 VSS A1 N_MM2_g N_A1_1 N_A1_6 N_A1_5 N_A1_8
+ PM_AO21x2_ASAP7_75t_R%A1
x_PM_AO21x2_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_AO21x2_ASAP7_75t_R%noxref_12
cc_28 N_noxref_12_1 N_MM7@2_g 0.00147148f
cc_29 N_noxref_12_1 N_Y_7 0.000494222f
x_PM_AO21x2_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_AO21x2_ASAP7_75t_R%noxref_13
cc_30 N_noxref_13_1 N_MM7@2_g 0.00147796f
cc_31 N_noxref_13_1 N_Y_8 0.00051415f
cc_32 N_noxref_13_1 N_noxref_12_1 0.00178634f
x_PM_AO21x2_ASAP7_75t_R%Y VSS Y N_MM7_d N_MM7@2_d N_MM8_d N_MM8@2_d N_Y_7 N_Y_9
+ N_Y_11 N_Y_2 N_Y_1 N_Y_12 N_Y_8 PM_AO21x2_ASAP7_75t_R%Y
cc_33 N_Y_7 N_NET16_16 0.000564264f
cc_34 N_Y_9 N_NET16_13 0.000870799f
cc_35 N_Y_11 N_NET16_1 0.00137431f
cc_36 N_Y_2 N_MM7@2_g 0.00223656f
cc_37 N_Y_9 N_NET16_17 0.00303559f
cc_38 N_Y_1 N_MM7@2_g 0.00304731f
cc_39 N_Y_12 N_NET16_15 0.00527859f
cc_40 N_Y_8 N_NET16_1 0.0054523f
cc_41 N_Y_8 N_MM7@2_g 0.0295456f
cc_42 N_Y_7 N_MM7_g 0.0367307f
cc_43 N_Y_7 N_MM7@2_g 0.0695411f
x_PM_AO21x2_ASAP7_75t_R%NET16 VSS N_MM7_g N_MM7@2_g N_MM3_d N_MM4_d N_MM1_s
+ N_MM5_s N_NET16_3 N_NET16_12 N_NET16_13 N_NET16_14 N_NET16_4 N_NET16_11
+ N_NET16_15 N_NET16_16 N_NET16_1 N_NET16_17 PM_AO21x2_ASAP7_75t_R%NET16
cc_44 N_NET16_3 N_A1_1 0.000398966f
cc_45 N_NET16_12 N_A1_1 0.000884153f
cc_46 N_NET16_3 N_MM2_g 0.000947351f
cc_47 N_NET16_13 N_A1_6 0.00125118f
cc_48 N_NET16_12 N_MM2_g 0.0362462f
cc_49 N_NET16_14 N_A2 0.000592474f
cc_50 N_NET16_3 N_A2_1 0.000592884f
cc_51 N_NET16_3 N_MM3_g 0.000918082f
cc_52 N_NET16_13 N_A2 0.00121539f
cc_53 N_NET16_12 N_A2_1 0.00144989f
cc_54 N_NET16_4 N_MM3_g 0.00160432f
cc_55 N_NET16_4 N_A2 0.00256596f
cc_56 N_NET16_12 N_MM3_g 0.015262f
cc_57 N_NET16_11 N_MM3_g 0.0550955f
cc_58 N_NET16_4 N_MM4_g 0.00198715f
cc_59 N_NET16_14 N_B_4 0.00107146f
cc_60 N_NET16_13 N_B_4 0.00123987f
cc_61 N_NET16_11 N_B_1 0.001259f
cc_62 N_MM7_g N_MM4_g 0.00163332f
cc_63 N_NET16_15 N_B_4 0.00616386f
cc_64 N_NET16_11 N_MM4_g 0.0374467f
*END of AO21x2_ASAP7_75t_R.pxi
.ENDS
** Design:	AO221x1_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AO221x1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AO221x1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AO221x1_ASAP7_75t_R%NET23 VSS 2 3 1
c1 1 VSS 0.00083422f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0540 $X2=0.1080 $Y2=0.0540
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0540 $X2=0.1080 $Y2=0.0540
.ends

.subckt PM_AO221x1_ASAP7_75t_R%NET24 VSS 2 3 1
c1 1 VSS 0.000837112f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0540 $X2=0.2700 $Y2=0.0540
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0540 $X2=0.2700 $Y2=0.0540
.ends

.subckt PM_AO221x1_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.0427062f
.ends

.subckt PM_AO221x1_ASAP7_75t_R%B2 VSS 6 3 1 4
c1 1 VSS 0.00556518f
c2 3 VSS 0.0353335f
c3 4 VSS 0.00429886f
r1 7 8 4.02252 $w=1.3e-08 $l=1.73e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1177 $X2=0.1350 $Y2=0.1350
r2 6 7 2.04041 $w=1.3e-08 $l=8.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1090 $X2=0.1350 $Y2=0.1177
r3 6 4 4.6055 $w=1.3e-08 $l=1.98e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1090 $X2=0.1350 $Y2=0.0892
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AO221x1_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00564971f
.ends

.subckt PM_AO221x1_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.0044513f
.ends

.subckt PM_AO221x1_ASAP7_75t_R%B1 VSS 8 3 1 4
c1 1 VSS 0.00603459f
c2 3 VSS 0.0081834f
c3 4 VSS 0.00386517f
r1 8 7 0.524677 $w=1.3e-08 $l=2.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1480 $X2=0.0810 $Y2=0.1457
r2 6 7 2.50679 $w=1.3e-08 $l=1.07e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1457
r3 4 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0980 $X2=0.0810 $Y2=0.1350
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r5 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AO221x1_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.00458339f
.ends

.subckt PM_AO221x1_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.00481978f
.ends

.subckt PM_AO221x1_ASAP7_75t_R%Y VSS 20 14 30 7 2 1 8 10
c1 1 VSS 0.00811434f
c2 2 VSS 0.00856484f
c3 7 VSS 0.00377533f
c4 8 VSS 0.00382743f
c5 9 VSS 0.00502436f
c6 10 VSS 0.00392983f
c7 11 VSS 0.00609556f
c8 12 VSS 0.00286209f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4840 $Y2=0.2025
r2 30 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r3 2 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2025
+ $X2=0.4860 $Y2=0.2340
r4 26 27 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.2340 $X2=0.4995 $Y2=0.2340
r5 11 24 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.2340 $X2=0.5130 $Y2=0.2160
r6 11 27 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.2340 $X2=0.4995 $Y2=0.2340
r7 23 24 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1980 $X2=0.5130 $Y2=0.2160
r8 22 23 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1765 $X2=0.5130 $Y2=0.1980
r9 21 22 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1560 $X2=0.5130 $Y2=0.1765
r10 20 21 1.98211 $w=1.3e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1475 $X2=0.5130 $Y2=0.1560
r11 20 19 0.46638 $w=1.3e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1475 $X2=0.5130 $Y2=0.1455
r12 18 19 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1455
r13 10 12 9.89378 $w=1.47818e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.0855 $X2=0.5130 $Y2=0.0360
r14 10 18 11.5429 $w=1.3e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0855 $X2=0.5130 $Y2=0.1350
r15 12 17 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.0360 $X2=0.4995 $Y2=0.0360
r16 16 17 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.0360 $X2=0.4995 $Y2=0.0360
r17 15 16 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4755
+ $Y=0.0360 $X2=0.4860 $Y2=0.0360
r18 9 15 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4665
+ $Y=0.0360 $X2=0.4755 $Y2=0.0360
r19 1 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0675
+ $X2=0.4860 $Y2=0.0360
r20 7 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0675 $X2=0.4840 $Y2=0.0675
r21 14 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4715 $Y2=0.0675
.ends

.subckt PM_AO221x1_ASAP7_75t_R%YN VSS 12 50 51 55 63 64 13 4 3 18 17 15 16 5 14
+ 24 19 22 20 23 1
c1 1 VSS 0.00428243f
c2 3 VSS 0.00568598f
c3 4 VSS 0.00298737f
c4 5 VSS 0.0074597f
c5 12 VSS 0.0805625f
c6 13 VSS 0.00329124f
c7 14 VSS 0.00403142f
c8 15 VSS 0.00305601f
c9 16 VSS 0.00375637f
c10 17 VSS 0.0345859f
c11 18 VSS 0.00108041f
c12 19 VSS 0.00422381f
c13 20 VSS 0.00230223f
c14 21 VSS 0.00306091f
c15 22 VSS 0.00111384f
c16 23 VSS 0.00310867f
c17 24 VSS 0.00173172f
r1 64 62 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r2 4 62 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r3 15 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r4 63 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
r5 4 59 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.1980
r6 58 59 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.1980 $X2=0.1080 $Y2=0.1980
r7 57 58 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1980 $X2=0.0945 $Y2=0.1980
r8 56 57 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.0555
+ $Y=0.1980 $X2=0.0810 $Y2=0.1980
r9 18 22 0.79938 $w=1.72857e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0375 $Y=0.1980 $X2=0.0270 $Y2=0.1980
r10 18 56 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0375
+ $Y=0.1980 $X2=0.0555 $Y2=0.1980
r11 22 53 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1980 $X2=0.0270 $Y2=0.1765
r12 55 54 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r13 13 54 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r14 52 53 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1170 $X2=0.0270 $Y2=0.1765
r15 16 21 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0575 $X2=0.0270 $Y2=0.0360
r16 16 52 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0575 $X2=0.0270 $Y2=0.1170
r17 51 49 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0540 $X2=0.2305 $Y2=0.0540
r18 5 49 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.0540 $X2=0.2305 $Y2=0.0540
r19 14 5 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0540 $X2=0.2160 $Y2=0.0540
r20 50 14 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0540 $X2=0.2015 $Y2=0.0540
r21 3 46 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0540 $Y2=0.0360
r22 21 45 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0360 $X2=0.0405 $Y2=0.0360
r23 5 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0540
+ $X2=0.2160 $Y2=0.0360
r24 46 47 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.0360 $X2=0.0675 $Y2=0.0360
r25 45 46 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r26 44 47 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0360 $X2=0.0675 $Y2=0.0360
r27 43 44 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.0810 $Y2=0.0360
r28 42 43 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1080 $Y2=0.0360
r29 41 42 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1600
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r30 40 41 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1780
+ $Y=0.0360 $X2=0.1600 $Y2=0.0360
r31 39 40 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.1780 $Y2=0.0360
r32 38 39 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1990
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r33 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.2295 $Y2=0.0360
r34 35 36 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2035
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r35 35 38 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2035
+ $Y=0.0360 $X2=0.1990 $Y2=0.0360
r36 34 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2295 $Y2=0.0360
r37 33 34 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r38 32 33 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r39 31 32 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3225
+ $Y=0.0360 $X2=0.2970 $Y2=0.0360
r40 17 23 7.0955 $w=1.42e-08 $l=3.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.3675
+ $Y=0.0360 $X2=0.4050 $Y2=0.0360
r41 17 31 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3675
+ $Y=0.0360 $X2=0.3225 $Y2=0.0360
r42 23 30 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.0360 $X2=0.4050 $Y2=0.0575
r43 19 24 6.97891 $w=1.53838e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.0980 $X2=0.4050 $Y2=0.1350
r44 19 30 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0980 $X2=0.4050 $Y2=0.0575
r45 20 26 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.1350 $X2=0.4545 $Y2=0.1350
r46 20 24 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4320 $Y=0.1350 $X2=0.4050 $Y2=0.1350
r47 12 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r48 1 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1350
+ $X2=0.4545 $Y2=0.1350
r49 3 13 1e-05
.ends

.subckt PM_AO221x1_ASAP7_75t_R%A1 VSS 8 3 1 4
c1 1 VSS 0.00670593f
c2 3 VSS 0.0456482f
c3 4 VSS 0.00367211f
r1 8 7 0.874462 $w=1.3e-08 $l=3.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1510 $X2=0.2430 $Y2=0.1472
r2 6 7 2.85657 $w=1.3e-08 $l=1.22e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1472
r3 4 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0980 $X2=0.2430 $Y2=0.1350
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r5 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AO221x1_ASAP7_75t_R%A2 VSS 6 3 1 4
c1 1 VSS 0.006277f
c2 3 VSS 0.072745f
c3 4 VSS 0.00427243f
r1 7 8 2.39019 $w=1.3e-08 $l=1.03e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1247 $X2=0.2970 $Y2=0.1350
r2 6 7 0.408082 $w=1.3e-08 $l=1.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1230 $X2=0.2970 $Y2=0.1247
r3 6 4 6.23783 $w=1.3e-08 $l=2.68e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1230 $X2=0.2970 $Y2=0.0962
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_AO221x1_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.00707858f
.ends

.subckt PM_AO221x1_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.0316643f
.ends

.subckt PM_AO221x1_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.0418102f
.ends

.subckt PM_AO221x1_ASAP7_75t_R%C VSS 6 3 1 4
c1 1 VSS 0.00662768f
c2 3 VSS 0.0347657f
c3 4 VSS 0.00450635f
r1 7 8 2.39019 $w=1.3e-08 $l=1.03e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1247 $X2=0.1890 $Y2=0.1350
r2 6 7 0.408082 $w=1.3e-08 $l=1.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1230 $X2=0.1890 $Y2=0.1247
r3 6 4 6.23783 $w=1.3e-08 $l=2.68e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1230 $X2=0.1890 $Y2=0.0962
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AO221x1_ASAP7_75t_R%S1 VSS 11 22 23 9 7 1 8 2
c1 1 VSS 0.00616531f
c2 2 VSS 0.00804606f
c3 7 VSS 0.00333233f
c4 8 VSS 0.0037193f
c5 9 VSS 0.00825084f
r1 23 21 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r2 1 21 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r3 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r4 22 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r5 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.1980
r6 18 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1980 $X2=0.2295 $Y2=0.1980
r7 16 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1980 $X2=0.2295 $Y2=0.1980
r8 15 16 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1980 $X2=0.2430 $Y2=0.1980
r9 14 15 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1980 $X2=0.2700 $Y2=0.1980
r10 9 12 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.3100
+ $Y=0.1980 $X2=0.3230 $Y2=0.1980
r11 9 14 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.3100
+ $Y=0.1980 $X2=0.2970 $Y2=0.1980
r12 2 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3230 $Y2=0.1980
r13 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3220 $Y2=0.2025
r14 11 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
.ends

.subckt PM_AO221x1_ASAP7_75t_R%S2 VSS 11 20 21 7 1 8 2 9
c1 1 VSS 0.00522071f
c2 2 VSS 0.00480622f
c3 7 VSS 0.00221667f
c4 8 VSS 0.00215959f
c5 9 VSS 0.0115194f
r1 21 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r2 2 19 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r4 20 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r5 2 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r6 15 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r7 14 15 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1485 $Y2=0.2340
r8 13 14 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r9 12 13 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2340 $X2=0.0945 $Y2=0.2340
r10 9 12 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0420
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r11 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r12 11 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r13 7 10 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r14 1 7 1e-05
.ends


*
.SUBCKT AO221x1_ASAP7_75t_R VSS VDD B1 B2 C A1 A2 Y
*
* VSS VSS
* VDD VDD
* B1 B1
* B2 B2
* C C
* A1 A1
* A2 A2
* Y Y
*
*

MM26 N_MM26_d N_MM26_g N_MM26_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM27 N_MM27_d N_MM27_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM28 N_MM28_d N_MM28_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2 N_MM2_d N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM0 N_MM0_d N_MM31_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM4 N_MM4_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM30 N_MM30_d N_MM26_g N_MM30_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM32 N_MM32_d N_MM27_g N_MM32_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM28_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM29 N_MM29_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM31 N_MM31_d N_MM31_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AO221x1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AO221x1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AO221x1_ASAP7_75t_R%NET23 VSS N_MM26_s N_MM27_d N_NET23_1
+ PM_AO221x1_ASAP7_75t_R%NET23
cc_1 N_NET23_1 N_MM26_g 0.0126336f
cc_2 N_NET23_1 N_MM27_g 0.012702f
x_PM_AO221x1_ASAP7_75t_R%NET24 VSS N_MM2_s N_MM0_d N_NET24_1
+ PM_AO221x1_ASAP7_75t_R%NET24
cc_3 N_NET24_1 N_MM2_g 0.0126402f
cc_4 N_NET24_1 N_MM31_g 0.0127119f
x_PM_AO221x1_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_AO221x1_ASAP7_75t_R%noxref_18
cc_5 N_noxref_18_1 N_MM3_g 0.00172066f
cc_6 N_noxref_18_1 N_noxref_16_1 0.00769805f
x_PM_AO221x1_ASAP7_75t_R%B2 VSS B2 N_MM27_g N_B2_1 N_B2_4
+ PM_AO221x1_ASAP7_75t_R%B2
cc_7 N_B2_1 N_B1_1 0.00130334f
cc_8 N_B2_4 N_B1_4 0.00354437f
cc_9 N_MM27_g N_MM26_g 0.00760991f
x_PM_AO221x1_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_AO221x1_ASAP7_75t_R%noxref_15
cc_10 N_noxref_15_1 N_MM26_g 0.00159575f
cc_11 N_noxref_15_1 N_YN_15 0.00088479f
cc_12 N_noxref_15_1 N_S2_7 0.0363593f
cc_13 N_noxref_15_1 N_noxref_14_1 0.00189854f
x_PM_AO221x1_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_AO221x1_ASAP7_75t_R%noxref_14
cc_14 N_noxref_14_1 N_MM26_g 0.00349958f
cc_15 N_noxref_14_1 N_YN_3 0.000436163f
cc_16 N_noxref_14_1 N_YN_13 0.0277832f
cc_17 N_noxref_14_1 N_S2_7 0.000581328f
x_PM_AO221x1_ASAP7_75t_R%B1 VSS B1 N_MM26_g N_B1_1 N_B1_4
+ PM_AO221x1_ASAP7_75t_R%B1
x_PM_AO221x1_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_AO221x1_ASAP7_75t_R%noxref_20
cc_18 N_noxref_20_1 N_MM3_g 0.00145273f
cc_19 N_noxref_20_1 N_Y_7 0.0385669f
x_PM_AO221x1_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_AO221x1_ASAP7_75t_R%noxref_21
cc_20 N_noxref_21_1 N_MM3_g 0.00145539f
cc_21 N_noxref_21_1 N_Y_8 0.0383939f
cc_22 N_noxref_21_1 N_noxref_20_1 0.00176866f
x_PM_AO221x1_ASAP7_75t_R%Y VSS Y N_MM4_d N_MM3_d N_Y_7 N_Y_2 N_Y_1 N_Y_8 N_Y_10
+ PM_AO221x1_ASAP7_75t_R%Y
cc_23 N_Y_7 N_YN_20 0.000190149f
cc_24 N_Y_7 N_YN_19 0.000651297f
cc_25 N_Y_7 N_YN_23 0.000778539f
cc_26 N_Y_2 N_MM3_g 0.00109815f
cc_27 N_Y_1 N_YN_1 0.00112703f
cc_28 N_Y_1 N_MM3_g 0.001168f
cc_29 N_Y_8 N_YN_1 0.00160963f
cc_30 N_Y_10 N_YN_20 0.00378296f
cc_31 N_Y_8 N_MM3_g 0.0152131f
cc_32 N_Y_7 N_MM3_g 0.054931f
x_PM_AO221x1_ASAP7_75t_R%YN VSS N_MM3_g N_MM28_d N_MM2_d N_MM26_d N_MM30_s
+ N_MM32_s N_YN_13 N_YN_4 N_YN_3 N_YN_18 N_YN_17 N_YN_15 N_YN_16 N_YN_5 N_YN_14
+ N_YN_24 N_YN_19 N_YN_22 N_YN_20 N_YN_23 N_YN_1 PM_AO221x1_ASAP7_75t_R%YN
cc_33 N_YN_13 N_MM26_g 0.0113736f
cc_34 N_YN_4 N_B1_1 0.000715597f
cc_35 N_YN_4 N_MM26_g 0.000907986f
cc_36 N_YN_3 N_MM26_g 0.000948084f
cc_37 N_YN_18 N_B1_4 0.00110783f
cc_38 N_YN_17 N_B1_4 0.00120711f
cc_39 N_YN_15 N_B1_1 0.00121304f
cc_40 N_YN_16 N_B1_4 0.00649649f
cc_41 N_YN_15 N_MM26_g 0.04915f
cc_42 N_YN_3 N_MM27_g 0.000192724f
cc_43 N_YN_4 N_MM27_g 0.00127552f
cc_44 N_YN_18 N_B2_4 0.000637692f
cc_45 N_YN_15 N_B2_1 0.000810704f
cc_46 N_YN_17 N_B2_4 0.00130846f
cc_47 N_YN_4 N_B2_4 0.00236286f
cc_48 N_YN_15 N_MM27_g 0.035528f
cc_49 N_YN_5 N_MM28_g 0.000660584f
cc_50 N_YN_17 N_C_4 0.00119644f
cc_51 N_YN_5 N_C_4 0.00169541f
cc_52 N_YN_14 N_MM28_g 0.0257642f
cc_53 N_YN_5 N_MM2_g 0.000939449f
cc_54 N_YN_17 N_A1_4 0.00130265f
cc_55 N_YN_5 N_A1_4 0.00169211f
cc_56 N_YN_14 N_MM2_g 0.0261987f
cc_57 N_YN_5 N_A2_4 0.000185407f
cc_58 N_YN_24 N_A2_4 0.000190458f
cc_59 N_YN_14 N_A2_4 0.000289686f
cc_60 N_YN_19 N_A2_4 0.000339916f
cc_61 N_YN_17 N_A2_4 0.00392866f
x_PM_AO221x1_ASAP7_75t_R%A1 VSS A1 N_MM2_g N_A1_1 N_A1_4
+ PM_AO221x1_ASAP7_75t_R%A1
cc_62 N_A1_1 N_C_1 0.00133605f
cc_63 N_A1_4 N_C_4 0.00345463f
cc_64 N_MM2_g N_MM28_g 0.00625088f
x_PM_AO221x1_ASAP7_75t_R%A2 VSS A2 N_MM31_g N_A2_1 N_A2_4
+ PM_AO221x1_ASAP7_75t_R%A2
cc_65 N_A2_1 N_A1_1 0.00145259f
cc_66 N_A2_4 N_A1_4 0.00336682f
cc_67 N_MM31_g N_MM2_g 0.00749733f
x_PM_AO221x1_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_AO221x1_ASAP7_75t_R%noxref_17
cc_68 N_noxref_17_1 N_MM31_g 0.00152859f
cc_69 N_noxref_17_1 N_S1_8 0.0357893f
cc_70 N_noxref_17_1 N_noxref_16_1 0.00135513f
x_PM_AO221x1_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_AO221x1_ASAP7_75t_R%noxref_16
cc_71 N_noxref_16_1 N_MM31_g 0.0034516f
cc_72 N_noxref_16_1 N_MM3_g 0.000504999f
cc_73 N_noxref_16_1 N_S1_8 0.000511078f
x_PM_AO221x1_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_AO221x1_ASAP7_75t_R%noxref_19
cc_74 N_noxref_19_1 N_MM3_g 0.00152922f
cc_75 N_noxref_19_1 N_S1_8 0.00061987f
cc_76 N_noxref_19_1 N_noxref_16_1 0.000472938f
cc_77 N_noxref_19_1 N_noxref_17_1 0.00766396f
cc_78 N_noxref_19_1 N_noxref_18_1 0.00123705f
x_PM_AO221x1_ASAP7_75t_R%C VSS C N_MM28_g N_C_1 N_C_4 PM_AO221x1_ASAP7_75t_R%C
cc_79 N_C_1 N_B2_1 0.0012141f
cc_80 N_C_4 N_B2_4 0.00350699f
cc_81 N_MM28_g N_MM27_g 0.0063593f
x_PM_AO221x1_ASAP7_75t_R%S1 VSS N_MM31_d N_MM1_d N_MM29_d N_S1_9 N_S1_7 N_S1_1
+ N_S1_8 N_S1_2 PM_AO221x1_ASAP7_75t_R%S1
cc_82 N_S1_9 N_MM28_g 0.00061811f
cc_83 N_S1_7 N_C_1 0.000801353f
cc_84 N_S1_1 N_C_4 0.000837787f
cc_85 N_S1_1 N_MM28_g 0.000881876f
cc_86 N_S1_7 N_MM28_g 0.0338891f
cc_87 N_S1_7 N_A1_1 0.000837116f
cc_88 N_S1_1 N_MM2_g 0.000883682f
cc_89 N_S1_9 N_A1_4 0.00114115f
cc_90 N_S1_1 N_A1_4 0.00128128f
cc_91 N_S1_7 N_MM2_g 0.0340191f
cc_92 N_S1_8 N_A2_1 0.000977683f
cc_93 N_S1_2 N_MM31_g 0.00108979f
cc_94 N_S1_9 N_A2_4 0.00129367f
cc_95 N_S1_2 N_A2_4 0.0015087f
cc_96 N_S1_8 N_MM31_g 0.0343348f
cc_97 N_S1_7 N_S2_8 0.000558588f
cc_98 N_S1_9 N_S2_9 0.00109636f
cc_99 N_S1_1 N_S2_2 0.00394044f
x_PM_AO221x1_ASAP7_75t_R%S2 VSS N_MM30_d N_MM32_d N_MM1_s N_S2_7 N_S2_1 N_S2_8
+ N_S2_2 N_S2_9 PM_AO221x1_ASAP7_75t_R%S2
cc_100 N_S2_7 N_B1_1 0.000725924f
cc_101 N_S2_1 N_MM26_g 0.00105932f
cc_102 N_S2_7 N_MM26_g 0.0345181f
cc_103 N_S2_8 N_B2_1 0.000662624f
cc_104 N_S2_2 N_MM27_g 0.000945592f
cc_105 N_S2_8 N_MM27_g 0.0346579f
cc_106 N_S2_8 N_C_1 0.000745827f
cc_107 N_S2_2 N_MM28_g 0.000947397f
cc_108 N_S2_8 N_MM28_g 0.0345036f
cc_109 N_S2_9 N_YN_4 0.000951408f
cc_110 N_S2_9 N_YN_15 0.00056429f
cc_111 N_S2_9 N_YN_22 0.000634145f
cc_112 N_S2_1 N_YN_18 0.000647747f
cc_113 N_S2_1 N_YN_16 0.000708385f
cc_114 N_S2_7 N_YN_15 0.00071357f
cc_115 N_S2_8 N_YN_15 0.00112456f
cc_116 N_S2_1 N_YN_4 0.00243187f
cc_117 N_S2_2 N_YN_4 0.00421426f
cc_118 N_S2_9 N_YN_18 0.00823397f
*END of AO221x1_ASAP7_75t_R.pxi
.ENDS
** Design:	AO221x2_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AO221x2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AO221x2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AO221x2_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.00712057f
.ends

.subckt PM_AO221x2_ASAP7_75t_R%NET23 VSS 2 3 1
c1 1 VSS 0.000833742f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0540 $X2=0.1080 $Y2=0.0540
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0540 $X2=0.1080 $Y2=0.0540
.ends

.subckt PM_AO221x2_ASAP7_75t_R%NET24 VSS 2 3 1
c1 1 VSS 0.000836959f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0540 $X2=0.2700 $Y2=0.0540
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0540 $X2=0.2700 $Y2=0.0540
.ends

.subckt PM_AO221x2_ASAP7_75t_R%S1 VSS 12 13 23 9 7 1 8 2
c1 1 VSS 0.00616375f
c2 2 VSS 0.00802821f
c3 7 VSS 0.00333082f
c4 8 VSS 0.00373983f
c5 9 VSS 0.00804093f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3220 $Y2=0.2025
r2 23 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r3 2 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3230 $Y2=0.1980
r4 19 20 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.3100
+ $Y=0.1980 $X2=0.3230 $Y2=0.1980
r5 18 19 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1980 $X2=0.3100 $Y2=0.1980
r6 17 18 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1980 $X2=0.2970 $Y2=0.1980
r7 16 17 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1980 $X2=0.2700 $Y2=0.1980
r8 15 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.1980 $X2=0.2430 $Y2=0.1980
r9 14 15 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1980 $X2=0.2295 $Y2=0.1980
r10 9 14 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2035
+ $Y=0.1980 $X2=0.2160 $Y2=0.1980
r11 1 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.1980
r12 12 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r13 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r14 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r15 13 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
.ends

.subckt PM_AO221x2_ASAP7_75t_R%A2 VSS 6 3 1 4
c1 1 VSS 0.00630493f
c2 3 VSS 0.0727329f
c3 4 VSS 0.00431355f
r1 7 8 2.39019 $w=1.3e-08 $l=1.03e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1247 $X2=0.2970 $Y2=0.1350
r2 6 7 0.408082 $w=1.3e-08 $l=1.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1230 $X2=0.2970 $Y2=0.1247
r3 6 4 6.23783 $w=1.3e-08 $l=2.68e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1230 $X2=0.2970 $Y2=0.0962
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_AO221x2_ASAP7_75t_R%B2 VSS 6 3 1 4
c1 1 VSS 0.00546737f
c2 3 VSS 0.0352844f
c3 4 VSS 0.00421658f
r1 7 8 4.02252 $w=1.3e-08 $l=1.73e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1177 $X2=0.1350 $Y2=0.1350
r2 6 7 2.04041 $w=1.3e-08 $l=8.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1090 $X2=0.1350 $Y2=0.1177
r3 6 4 4.6055 $w=1.3e-08 $l=1.98e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1090 $X2=0.1350 $Y2=0.0892
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AO221x2_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.0427f
.ends

.subckt PM_AO221x2_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00565096f
.ends

.subckt PM_AO221x2_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.031667f
.ends

.subckt PM_AO221x2_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00445385f
.ends

.subckt PM_AO221x2_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.0418075f
.ends

.subckt PM_AO221x2_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.0425967f
.ends

.subckt PM_AO221x2_ASAP7_75t_R%A1 VSS 8 3 1 4
c1 1 VSS 0.00651904f
c2 3 VSS 0.0455577f
c3 4 VSS 0.00352515f
r1 8 7 0.874462 $w=1.3e-08 $l=3.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1510 $X2=0.2430 $Y2=0.1472
r2 6 7 2.85657 $w=1.3e-08 $l=1.22e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1472
r3 4 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0980 $X2=0.2430 $Y2=0.1350
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r5 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AO221x2_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.04259f
.ends

.subckt PM_AO221x2_ASAP7_75t_R%Y VSS 23 16 17 33 34 7 8 9 1 11 2
c1 1 VSS 0.00993714f
c2 2 VSS 0.0104584f
c3 7 VSS 0.00451893f
c4 8 VSS 0.00454916f
c5 9 VSS 0.00715504f
c6 10 VSS 0.00629323f
c7 11 VSS 0.00834241f
c8 12 VSS 0.00341781f
c9 13 VSS 0.00339498f
r1 34 32 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r2 2 32 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4860 $Y2=0.2025
r4 33 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r5 2 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2025
+ $X2=0.4860 $Y2=0.2340
r6 28 29 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.2340 $X2=0.5130 $Y2=0.2340
r7 10 28 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4755
+ $Y=0.2340 $X2=0.4860 $Y2=0.2340
r8 13 27 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.2340 $X2=0.5400 $Y2=0.2160
r9 13 29 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5400 $Y=0.2340 $X2=0.5130 $Y2=0.2340
r10 26 27 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1980 $X2=0.5400 $Y2=0.2160
r11 25 26 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1765 $X2=0.5400 $Y2=0.1980
r12 24 25 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1560 $X2=0.5400 $Y2=0.1765
r13 23 24 1.98211 $w=1.3e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1475 $X2=0.5400 $Y2=0.1560
r14 23 22 0.46638 $w=1.3e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1475 $X2=0.5400 $Y2=0.1455
r15 21 22 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1350 $X2=0.5400 $Y2=0.1455
r16 11 12 9.89378 $w=1.47818e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5400 $Y=0.0855 $X2=0.5400 $Y2=0.0360
r17 11 21 11.5429 $w=1.3e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.0855 $X2=0.5400 $Y2=0.1350
r18 12 20 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5400 $Y=0.0360 $X2=0.5130 $Y2=0.0360
r19 19 20 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.0360 $X2=0.5130 $Y2=0.0360
r20 18 19 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4755
+ $Y=0.0360 $X2=0.4860 $Y2=0.0360
r21 9 18 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4665
+ $Y=0.0360 $X2=0.4755 $Y2=0.0360
r22 1 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0675
+ $X2=0.4860 $Y2=0.0360
r23 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0675 $X2=0.5005 $Y2=0.0675
r24 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.0675 $X2=0.5005 $Y2=0.0675
r25 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0675 $X2=0.4860 $Y2=0.0675
r26 16 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4715 $Y2=0.0675
.ends

.subckt PM_AO221x2_ASAP7_75t_R%C VSS 6 3 1 4
c1 1 VSS 0.0066981f
c2 3 VSS 0.03481f
c3 4 VSS 0.00456067f
r1 7 8 2.39019 $w=1.3e-08 $l=1.03e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1247 $X2=0.1890 $Y2=0.1350
r2 6 7 0.408082 $w=1.3e-08 $l=1.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1230 $X2=0.1890 $Y2=0.1247
r3 6 4 6.23783 $w=1.3e-08 $l=2.68e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1230 $X2=0.1890 $Y2=0.0962
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AO221x2_ASAP7_75t_R%B1 VSS 8 3 1 4
c1 1 VSS 0.0060299f
c2 3 VSS 0.00818105f
c3 4 VSS 0.00384377f
r1 8 7 0.524677 $w=1.3e-08 $l=2.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1480 $X2=0.0810 $Y2=0.1457
r2 6 7 2.50679 $w=1.3e-08 $l=1.07e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1457
r3 4 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0980 $X2=0.0810 $Y2=0.1350
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r5 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AO221x2_ASAP7_75t_R%S2 VSS 11 20 21 7 1 8 2 9
c1 1 VSS 0.00522271f
c2 2 VSS 0.00480395f
c3 7 VSS 0.00221886f
c4 8 VSS 0.00216168f
c5 9 VSS 0.0115304f
r1 21 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r2 2 19 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r4 20 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r5 2 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r6 15 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r7 14 15 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1485 $Y2=0.2340
r8 13 14 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r9 12 13 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2340 $X2=0.0945 $Y2=0.2340
r10 9 12 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0420
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r11 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r12 11 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r13 7 10 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r14 1 7 1e-05
.ends

.subckt PM_AO221x2_ASAP7_75t_R%YN VSS 12 13 61 62 66 74 75 14 4 3 19 16 18 17 5
+ 15 25 20 23 21 1 24
c1 1 VSS 0.00847902f
c2 3 VSS 0.00595184f
c3 4 VSS 0.0030101f
c4 5 VSS 0.00748942f
c5 12 VSS 0.0813045f
c6 13 VSS 0.0807074f
c7 14 VSS 0.00457739f
c8 15 VSS 0.00525537f
c9 16 VSS 0.00464782f
c10 17 VSS 0.00627287f
c11 18 VSS 0.036474f
c12 19 VSS 0.00158709f
c13 20 VSS 0.00477312f
c14 21 VSS 0.00308866f
c15 22 VSS 0.00349456f
c16 23 VSS 0.00168012f
c17 24 VSS 0.00332277f
c18 25 VSS 0.00190641f
r1 75 73 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r2 4 73 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r3 16 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r4 74 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
r5 4 70 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.1980
r6 69 70 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.1980 $X2=0.1080 $Y2=0.1980
r7 68 69 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1980 $X2=0.0945 $Y2=0.1980
r8 67 68 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.0555
+ $Y=0.1980 $X2=0.0810 $Y2=0.1980
r9 19 23 0.79938 $w=1.72857e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0375 $Y=0.1980 $X2=0.0270 $Y2=0.1980
r10 19 67 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0375
+ $Y=0.1980 $X2=0.0555 $Y2=0.1980
r11 23 64 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1980 $X2=0.0270 $Y2=0.1765
r12 66 65 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r13 14 65 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r14 63 64 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1170 $X2=0.0270 $Y2=0.1765
r15 17 22 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0575 $X2=0.0270 $Y2=0.0360
r16 17 63 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0575 $X2=0.0270 $Y2=0.1170
r17 62 60 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0540 $X2=0.2305 $Y2=0.0540
r18 5 60 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.0540 $X2=0.2305 $Y2=0.0540
r19 15 5 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0540 $X2=0.2160 $Y2=0.0540
r20 61 15 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0540 $X2=0.2015 $Y2=0.0540
r21 3 57 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0540 $Y2=0.0360
r22 22 56 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0360 $X2=0.0405 $Y2=0.0360
r23 5 47 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0540
+ $X2=0.2160 $Y2=0.0360
r24 57 58 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.0360 $X2=0.0675 $Y2=0.0360
r25 56 57 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r26 55 58 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0360 $X2=0.0675 $Y2=0.0360
r27 54 55 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.0810 $Y2=0.0360
r28 53 54 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1080 $Y2=0.0360
r29 52 53 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1600
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r30 51 52 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1780
+ $Y=0.0360 $X2=0.1600 $Y2=0.0360
r31 50 51 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.1780 $Y2=0.0360
r32 49 50 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1990
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r33 47 48 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.2295 $Y2=0.0360
r34 46 47 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2035
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r35 46 49 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2035
+ $Y=0.0360 $X2=0.1990 $Y2=0.0360
r36 45 48 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2295 $Y2=0.0360
r37 44 45 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r38 43 44 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r39 42 43 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3225
+ $Y=0.0360 $X2=0.2970 $Y2=0.0360
r40 18 24 7.0955 $w=1.42e-08 $l=3.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.3675
+ $Y=0.0360 $X2=0.4050 $Y2=0.0360
r41 18 42 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3675
+ $Y=0.0360 $X2=0.3225 $Y2=0.0360
r42 24 41 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.0360 $X2=0.4050 $Y2=0.0575
r43 20 25 6.97891 $w=1.53838e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.0980 $X2=0.4050 $Y2=0.1350
r44 20 41 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0980 $X2=0.4050 $Y2=0.0575
r45 13 34 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r46 21 36 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.1350 $X2=0.4545 $Y2=0.1350
r47 21 25 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4320 $Y=0.1350 $X2=0.4050 $Y2=0.1350
r48 32 34 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5005 $Y=0.1350 $X2=0.5130 $Y2=0.1350
r49 31 32 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4860 $Y=0.1350 $X2=0.5005 $Y2=0.1350
r50 30 31 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4715 $Y=0.1350 $X2=0.4860 $Y2=0.1350
r51 28 30 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.4685 $Y=0.1350 $X2=0.4715 $Y2=0.1350
r52 27 28 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4685 $Y2=0.1350
r53 27 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1350
+ $X2=0.4545 $Y2=0.1350
r54 1 27 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.4495
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r55 1 29 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.4495
+ $Y=0.1350 $X2=0.4485 $Y2=0.1350
r56 12 27 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4590 $Y2=0.1350
r57 12 29 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.4590 $Y=0.1350 $X2=0.4485 $Y2=0.1350
r58 12 30 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4715 $Y2=0.1350
r59 3 14 1e-05
.ends


*
.SUBCKT AO221x2_ASAP7_75t_R VSS VDD B1 B2 C A1 A2 Y
*
* VSS VSS
* VDD VDD
* B1 B1
* B2 B2
* C C
* A1 A1
* A2 A2
* Y Y
*
*

MM26 N_MM26_d N_MM26_g N_MM26_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM27 N_MM27_d N_MM27_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM28 N_MM28_d N_MM28_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2 N_MM2_d N_MM29_g N_MM2_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM0 N_MM0_d N_MM31_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM4 N_MM4_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@2 N_MM4@2_d N_MM3@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM30 N_MM30_d N_MM26_g N_MM30_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM32 N_MM32_d N_MM27_g N_MM32_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM28_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM29 N_MM29_d N_MM29_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM31 N_MM31_d N_MM31_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3@2 N_MM3@2_d N_MM3@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AO221x2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AO221x2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AO221x2_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_AO221x2_ASAP7_75t_R%noxref_17
cc_1 N_noxref_17_1 N_MM31_g 0.00152868f
cc_2 N_noxref_17_1 N_S1_8 0.0357463f
cc_3 N_noxref_17_1 N_noxref_16_1 0.00134897f
x_PM_AO221x2_ASAP7_75t_R%NET23 VSS N_MM26_s N_MM27_d N_NET23_1
+ PM_AO221x2_ASAP7_75t_R%NET23
cc_4 N_NET23_1 N_MM26_g 0.0126216f
cc_5 N_NET23_1 N_MM27_g 0.0127144f
x_PM_AO221x2_ASAP7_75t_R%NET24 VSS N_MM2_s N_MM0_d N_NET24_1
+ PM_AO221x2_ASAP7_75t_R%NET24
cc_6 N_NET24_1 N_MM29_g 0.0126399f
cc_7 N_NET24_1 N_MM31_g 0.0127123f
x_PM_AO221x2_ASAP7_75t_R%S1 VSS N_MM29_d N_MM1_d N_MM31_d N_S1_9 N_S1_7 N_S1_1
+ N_S1_8 N_S1_2 PM_AO221x2_ASAP7_75t_R%S1
cc_8 N_S1_9 N_MM28_g 0.000601396f
cc_9 N_S1_7 N_C_1 0.000800989f
cc_10 N_S1_1 N_C_4 0.000837834f
cc_11 N_S1_1 N_MM28_g 0.000881476f
cc_12 N_S1_7 N_MM28_g 0.0338737f
cc_13 N_S1_7 N_A1_1 0.000836764f
cc_14 N_S1_1 N_MM29_g 0.000883281f
cc_15 N_S1_9 N_A1_4 0.00114466f
cc_16 N_S1_1 N_A1_4 0.0012358f
cc_17 N_S1_7 N_MM29_g 0.034003f
cc_18 N_S1_8 N_A2_1 0.000977239f
cc_19 N_S1_2 N_MM31_g 0.00108792f
cc_20 N_S1_9 N_A2_4 0.00128756f
cc_21 N_S1_2 N_A2_4 0.00152176f
cc_22 N_S1_8 N_MM31_g 0.0343133f
cc_23 N_S1_7 N_S2_8 0.000558334f
cc_24 N_S1_9 N_S2_9 0.00105023f
cc_25 N_S1_1 N_S2_2 0.00393865f
x_PM_AO221x2_ASAP7_75t_R%A2 VSS A2 N_MM31_g N_A2_1 N_A2_4
+ PM_AO221x2_ASAP7_75t_R%A2
cc_26 N_A2_1 N_A1_1 0.00145259f
cc_27 N_A2_4 N_A1_4 0.00341289f
cc_28 N_MM31_g N_MM29_g 0.00749733f
x_PM_AO221x2_ASAP7_75t_R%B2 VSS B2 N_MM27_g N_B2_1 N_B2_4
+ PM_AO221x2_ASAP7_75t_R%B2
cc_29 N_B2_1 N_B1_1 0.00130334f
cc_30 N_B2_4 N_B1_4 0.00351461f
cc_31 N_MM27_g N_MM26_g 0.00760991f
x_PM_AO221x2_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_AO221x2_ASAP7_75t_R%noxref_18
cc_32 N_noxref_18_1 N_MM3_g 0.00175675f
cc_33 N_noxref_18_1 N_noxref_16_1 0.00770153f
x_PM_AO221x2_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_AO221x2_ASAP7_75t_R%noxref_15
cc_34 N_noxref_15_1 N_MM26_g 0.00159547f
cc_35 N_noxref_15_1 N_YN_16 0.000878108f
cc_36 N_noxref_15_1 N_S2_7 0.0363703f
cc_37 N_noxref_15_1 N_noxref_14_1 0.00189586f
x_PM_AO221x2_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_AO221x2_ASAP7_75t_R%noxref_16
cc_38 N_noxref_16_1 N_MM31_g 0.00346014f
cc_39 N_noxref_16_1 N_MM3_g 0.000513831f
cc_40 N_noxref_16_1 N_S1_8 0.00050882f
x_PM_AO221x2_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_AO221x2_ASAP7_75t_R%noxref_14
cc_41 N_noxref_14_1 N_MM26_g 0.00349615f
cc_42 N_noxref_14_1 N_YN_17 0.000348236f
cc_43 N_noxref_14_1 N_YN_3 0.000436163f
cc_44 N_noxref_14_1 N_YN_14 0.0274093f
cc_45 N_noxref_14_1 N_S2_7 0.000580101f
x_PM_AO221x2_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_AO221x2_ASAP7_75t_R%noxref_19
cc_46 N_noxref_19_1 N_MM3_g 0.00155906f
cc_47 N_noxref_19_1 N_S1_8 0.000615876f
cc_48 N_noxref_19_1 N_noxref_16_1 0.000470823f
cc_49 N_noxref_19_1 N_noxref_17_1 0.0076588f
cc_50 N_noxref_19_1 N_noxref_18_1 0.00123888f
x_PM_AO221x2_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_AO221x2_ASAP7_75t_R%noxref_21
cc_51 N_noxref_21_1 N_MM3@2_g 0.00147435f
cc_52 N_noxref_21_1 N_Y_8 0.000530177f
cc_53 N_noxref_21_1 N_noxref_20_1 0.00178828f
x_PM_AO221x2_ASAP7_75t_R%A1 VSS A1 N_MM29_g N_A1_1 N_A1_4
+ PM_AO221x2_ASAP7_75t_R%A1
cc_54 N_A1_1 N_C_1 0.00133605f
cc_55 N_A1_4 N_C_4 0.00327267f
cc_56 N_MM29_g N_MM28_g 0.00625088f
x_PM_AO221x2_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_AO221x2_ASAP7_75t_R%noxref_20
cc_57 N_noxref_20_1 N_MM3@2_g 0.00148192f
cc_58 N_noxref_20_1 N_Y_7 0.000528348f
x_PM_AO221x2_ASAP7_75t_R%Y VSS Y N_MM4_d N_MM4@2_d N_MM3_d N_MM3@2_d N_Y_7
+ N_Y_8 N_Y_9 N_Y_1 N_Y_11 N_Y_2 PM_AO221x2_ASAP7_75t_R%Y
cc_59 N_Y_7 N_YN_25 0.000149656f
cc_60 N_Y_7 N_YN_21 0.000271745f
cc_61 N_Y_7 N_YN_20 0.000602307f
cc_62 N_Y_7 N_YN_1 0.000778716f
cc_63 N_Y_8 N_MM3@2_g 0.0305425f
cc_64 N_Y_9 N_YN_24 0.000880878f
cc_65 N_Y_1 N_YN_21 0.00128352f
cc_66 N_Y_11 N_YN_1 0.00147924f
cc_67 N_Y_2 N_MM3@2_g 0.00199991f
cc_68 N_Y_1 N_MM3@2_g 0.00207233f
cc_69 N_Y_8 N_YN_1 0.00480454f
cc_70 N_Y_7 N_MM3_g 0.0368593f
cc_71 N_Y_7 N_MM3@2_g 0.0676653f
x_PM_AO221x2_ASAP7_75t_R%C VSS C N_MM28_g N_C_1 N_C_4 PM_AO221x2_ASAP7_75t_R%C
cc_72 N_C_1 N_B2_1 0.0012141f
cc_73 N_C_4 N_B2_4 0.00347029f
cc_74 N_MM28_g N_MM27_g 0.0063593f
x_PM_AO221x2_ASAP7_75t_R%B1 VSS B1 N_MM26_g N_B1_1 N_B1_4
+ PM_AO221x2_ASAP7_75t_R%B1
x_PM_AO221x2_ASAP7_75t_R%S2 VSS N_MM30_d N_MM32_d N_MM1_s N_S2_7 N_S2_1 N_S2_8
+ N_S2_2 N_S2_9 PM_AO221x2_ASAP7_75t_R%S2
cc_75 N_S2_7 N_B1_1 0.000726156f
cc_76 N_S2_1 N_MM26_g 0.00105966f
cc_77 N_S2_7 N_MM26_g 0.0345298f
cc_78 N_S2_8 N_B2_1 0.000662835f
cc_79 N_S2_2 N_MM27_g 0.000945894f
cc_80 N_S2_8 N_MM27_g 0.0346633f
cc_81 N_S2_8 N_C_1 0.000746065f
cc_82 N_S2_2 N_MM28_g 0.0009477f
cc_83 N_S2_8 N_MM28_g 0.0345145f
cc_84 N_S2_9 N_YN_4 0.000951711f
cc_85 N_S2_9 N_YN_16 0.00056447f
cc_86 N_S2_9 N_YN_23 0.000633157f
cc_87 N_S2_1 N_YN_19 0.000647954f
cc_88 N_S2_1 N_YN_17 0.000699328f
cc_89 N_S2_7 N_YN_16 0.000713798f
cc_90 N_S2_8 N_YN_16 0.00112491f
cc_91 N_S2_1 N_YN_4 0.00243264f
cc_92 N_S2_2 N_YN_4 0.0042156f
cc_93 N_S2_9 N_YN_19 0.00823427f
x_PM_AO221x2_ASAP7_75t_R%YN VSS N_MM3_g N_MM3@2_g N_MM28_d N_MM2_d N_MM26_d
+ N_MM30_s N_MM32_s N_YN_14 N_YN_4 N_YN_3 N_YN_19 N_YN_16 N_YN_18 N_YN_17
+ N_YN_5 N_YN_15 N_YN_25 N_YN_20 N_YN_23 N_YN_21 N_YN_1 N_YN_24
+ PM_AO221x2_ASAP7_75t_R%YN
cc_94 N_YN_14 N_MM26_g 0.0113736f
cc_95 N_YN_4 N_B1_1 0.000715597f
cc_96 N_YN_4 N_MM26_g 0.000907986f
cc_97 N_YN_3 N_MM26_g 0.000948084f
cc_98 N_YN_19 N_B1_4 0.00110782f
cc_99 N_YN_16 N_B1_1 0.00121304f
cc_100 N_YN_18 N_B1_4 0.00127699f
cc_101 N_YN_17 N_B1_4 0.00663389f
cc_102 N_YN_16 N_MM26_g 0.0491509f
cc_103 N_YN_4 N_MM27_g 0.00143947f
cc_104 N_YN_3 N_MM27_g 0.000192724f
cc_105 N_YN_19 N_B2_4 0.00063767f
cc_106 N_YN_16 N_B2_1 0.000810704f
cc_107 N_YN_18 N_B2_4 0.00137761f
cc_108 N_YN_4 N_B2_4 0.00230462f
cc_109 N_YN_16 N_MM27_g 0.035366f
cc_110 N_YN_5 N_MM28_g 0.000804701f
cc_111 N_YN_18 N_C_4 0.00125793f
cc_112 N_YN_5 N_C_4 0.00170301f
cc_113 N_YN_15 N_MM28_g 0.0256217f
cc_114 N_YN_5 N_MM29_g 0.000939449f
cc_115 N_YN_18 N_A1_4 0.00135305f
cc_116 N_YN_5 N_A1_4 0.00163355f
cc_117 N_YN_15 N_MM29_g 0.0262104f
cc_118 N_YN_15 N_A2_4 0.000461147f
cc_119 N_YN_25 N_A2_4 0.000178198f
cc_120 N_YN_5 N_A2_4 0.000185407f
cc_121 N_YN_20 N_A2_4 0.000336542f
cc_122 N_YN_18 N_A2_4 0.00393322f
*END of AO221x2_ASAP7_75t_R.pxi
.ENDS
** Design:	AO222x2_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AO222x2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AO222x2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AO222x2_ASAP7_75t_R%NET36 VSS 2 3 1
c1 1 VSS 0.00101578f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_AO222x2_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.0430302f
.ends

.subckt PM_AO222x2_ASAP7_75t_R%NET37 VSS 2 3 1
c1 1 VSS 0.00101327f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2160 $Y2=0.0675
.ends

.subckt PM_AO222x2_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.00737871f
.ends

.subckt PM_AO222x2_ASAP7_75t_R%NET38 VSS 2 3 1
c1 1 VSS 0.00101358f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4320 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4320 $Y2=0.0675
.ends

.subckt PM_AO222x2_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.0423816f
.ends

.subckt PM_AO222x2_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.0047385f
.ends

.subckt PM_AO222x2_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.0423842f
.ends

.subckt PM_AO222x2_ASAP7_75t_R%Y VSS 26 18 19 34 35 7 8 12 13 10 2 1
c1 1 VSS 0.00873701f
c2 2 VSS 0.0106333f
c3 7 VSS 0.00454923f
c4 8 VSS 0.00456696f
c5 9 VSS 0.00982936f
c6 10 VSS 0.00139396f
c7 11 VSS 0.00661474f
c8 12 VSS 0.00747505f
c9 13 VSS 0.00256277f
c10 14 VSS 0.00346759f
c11 15 VSS 0.00349839f
r1 35 33 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r2 2 33 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5400 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.2025 $X2=0.5400 $Y2=0.2025
r4 34 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.2025 $X2=0.5255 $Y2=0.2025
r5 2 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.2025
+ $X2=0.5400 $Y2=0.2340
r6 30 31 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.2340 $X2=0.5515 $Y2=0.2340
r7 9 15 7.2121 $w=1.41842e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5830
+ $Y=0.2340 $X2=0.6210 $Y2=0.2340
r8 9 31 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5830
+ $Y=0.2340 $X2=0.5515 $Y2=0.2340
r9 15 28 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.2340 $X2=0.6210 $Y2=0.2125
r10 27 28 9.0361 $w=1.3e-08 $l=3.88e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1737 $X2=0.6210 $Y2=0.2125
r11 26 27 6.23783 $w=1.3e-08 $l=2.67e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1470 $X2=0.6210 $Y2=0.1737
r12 26 25 0.408082 $w=1.3e-08 $l=1.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1470 $X2=0.6210 $Y2=0.1452
r13 24 25 2.3902 $w=1.3e-08 $l=1.02e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1452
r14 23 24 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1035 $X2=0.6210 $Y2=0.1350
r15 12 14 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.0630 $X2=0.6210 $Y2=0.0360
r16 12 23 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0630 $X2=0.6210 $Y2=0.1035
r17 14 22 7.2121 $w=1.41842e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.0360 $X2=0.5830 $Y2=0.0360
r18 11 13 1.03257 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5515 $Y=0.0360 $X2=0.5400 $Y2=0.0360
r19 11 22 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5515
+ $Y=0.0360 $X2=0.5830 $Y2=0.0360
r20 10 20 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.0490 $X2=0.5400 $Y2=0.0620
r21 10 13 1.38235 $w=1.97846e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5400 $Y=0.0490 $X2=0.5400 $Y2=0.0360
r22 1 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.0675
+ $X2=0.5400 $Y2=0.0620
r23 19 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.0675 $X2=0.5545 $Y2=0.0675
r24 1 17 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5400 $Y=0.0675 $X2=0.5545 $Y2=0.0675
r25 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.0675 $X2=0.5400 $Y2=0.0675
r26 18 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.0675 $X2=0.5255 $Y2=0.0675
.ends

.subckt PM_AO222x2_ASAP7_75t_R%C2 VSS 8 3 1 4
c1 1 VSS 0.00663738f
c2 3 VSS 0.0461779f
c3 4 VSS 0.00448496f
r1 8 7 0.408082 $w=1.3e-08 $l=1.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1470 $X2=0.1350 $Y2=0.1452
r2 6 7 2.39019 $w=1.3e-08 $l=1.02e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1452
r3 4 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0980 $X2=0.1350 $Y2=0.1350
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r5 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AO222x2_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.00523242f
.ends

.subckt PM_AO222x2_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.00586705f
.ends

.subckt PM_AO222x2_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.00548473f
.ends

.subckt PM_AO222x2_ASAP7_75t_R%C1 VSS 6 3 1 4
c1 1 VSS 0.00724309f
c2 3 VSS 0.00881257f
c3 4 VSS 0.00455757f
r1 7 8 5.42166 $w=1.3e-08 $l=2.33e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1117 $X2=0.0810 $Y2=0.1350
r2 6 7 3.43955 $w=1.3e-08 $l=1.47e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0970 $X2=0.0810 $Y2=0.1117
r3 6 4 3.20636 $w=1.3e-08 $l=1.38e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0970 $X2=0.0810 $Y2=0.0832
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AO222x2_ASAP7_75t_R%NET23 VSS 15 16 66 68 72 80 81 20 3 4 23 22 21
+ 17 18 5 6 19 25 1 24 29 27 28
c1 1 VSS 0.00728007f
c2 3 VSS 0.00599286f
c3 4 VSS 0.00302884f
c4 5 VSS 0.00634179f
c5 6 VSS 0.00627876f
c6 15 VSS 0.080634f
c7 16 VSS 0.0808019f
c8 17 VSS 0.00417237f
c9 18 VSS 0.00445433f
c10 19 VSS 0.00474346f
c11 20 VSS 0.00357807f
c12 21 VSS 0.00453721f
c13 22 VSS 0.0425436f
c14 23 VSS 0.00150457f
c15 24 VSS 0.00250871f
c16 25 VSS 0.00144172f
c17 26 VSS 0.00309406f
c18 27 VSS 0.00131822f
c19 28 VSS 0.00279477f
c20 29 VSS 0.000507108f
r1 81 79 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r2 4 79 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r3 20 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r4 80 20 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
r5 4 76 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.1980
r6 75 76 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.1980 $X2=0.1080 $Y2=0.1980
r7 74 75 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1980 $X2=0.0945 $Y2=0.1980
r8 73 74 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.0560
+ $Y=0.1980 $X2=0.0810 $Y2=0.1980
r9 23 27 1.96533 $w=1.59032e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0335 $Y=0.1980 $X2=0.0180 $Y2=0.1980
r10 23 73 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0335
+ $Y=0.1980 $X2=0.0560 $Y2=0.1980
r11 27 70 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.1980 $X2=0.0180 $Y2=0.1765
r12 72 71 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r13 17 71 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r14 69 70 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1170 $X2=0.0180 $Y2=0.1765
r15 21 26 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.0575 $X2=0.0180 $Y2=0.0360
r16 21 69 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0575 $X2=0.0180 $Y2=0.1170
r17 18 5 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2680 $Y2=0.0675
r18 68 18 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
r19 66 65 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r20 19 65 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3800 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r21 3 63 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0540 $Y2=0.0360
r22 26 62 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0360 $X2=0.0360 $Y2=0.0360
r23 5 51 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2700 $Y2=0.0360
r24 6 48 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.0675
+ $X2=0.3780 $Y2=0.0360
r25 63 64 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.0360 $X2=0.0675 $Y2=0.0360
r26 62 63 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r27 61 64 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0360 $X2=0.0675 $Y2=0.0360
r28 60 61 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1060
+ $Y=0.0360 $X2=0.0810 $Y2=0.0360
r29 59 60 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1240
+ $Y=0.0360 $X2=0.1060 $Y2=0.0360
r30 58 59 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1240 $Y2=0.0360
r31 57 58 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r32 56 57 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r33 55 56 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2000
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r34 54 55 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2180
+ $Y=0.0360 $X2=0.2000 $Y2=0.0360
r35 53 54 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2180 $Y2=0.0360
r36 51 52 11.5429 $w=1.3e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.3195 $Y2=0.0360
r37 50 51 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r38 50 53 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r39 48 49 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0360 $X2=0.3915 $Y2=0.0360
r40 47 48 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3645
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r41 47 52 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3645
+ $Y=0.0360 $X2=0.3195 $Y2=0.0360
r42 46 49 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0360 $X2=0.3915 $Y2=0.0360
r43 45 46 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4050 $Y2=0.0360
r44 44 45 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r45 22 28 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4770
+ $Y=0.0360 $X2=0.4950 $Y2=0.0360
r46 22 44 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4770
+ $Y=0.0360 $X2=0.4590 $Y2=0.0360
r47 28 43 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4950 $Y=0.0360 $X2=0.4950 $Y2=0.0575
r48 42 43 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4950
+ $Y=0.0755 $X2=0.4950 $Y2=0.0575
r49 24 29 5.69636 $w=1.58e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4950 $Y=0.1035 $X2=0.4950 $Y2=0.1350
r50 24 42 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4950
+ $Y=0.1035 $X2=0.4950 $Y2=0.0755
r51 29 39 3.01468 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4950
+ $Y=0.1350 $X2=0.5150 $Y2=0.1350
r52 16 36 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1350
r53 38 39 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5285
+ $Y=0.1350 $X2=0.5150 $Y2=0.1350
r54 25 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5400 $Y=0.1350
+ $X2=0.5400 $Y2=0.1350
r55 25 38 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1350 $X2=0.5285 $Y2=0.1350
r56 34 36 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5545 $Y=0.1350 $X2=0.5670 $Y2=0.1350
r57 33 34 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5400 $Y=0.1350 $X2=0.5545 $Y2=0.1350
r58 32 33 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5255 $Y=0.1350 $X2=0.5400 $Y2=0.1350
r59 15 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r60 1 31 2.90696 $w=2.1681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5025 $Y2=0.1350
r61 1 32 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5255 $Y2=0.1350
r62 15 31 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.5130 $Y=0.1350 $X2=0.5025 $Y2=0.1350
r63 15 32 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5255 $Y2=0.1350
r64 3 17 1e-05
r65 6 19 1e-05
.ends

.subckt PM_AO222x2_ASAP7_75t_R%B1 VSS 8 3 1 4
c1 1 VSS 0.00775396f
c2 3 VSS 0.00932883f
c3 4 VSS 0.00520202f
r1 8 7 0.408082 $w=1.3e-08 $l=1.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1470 $X2=0.2430 $Y2=0.1452
r2 6 7 2.39019 $w=1.3e-08 $l=1.02e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1452
r3 4 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0980 $X2=0.2430 $Y2=0.1350
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r5 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AO222x2_ASAP7_75t_R%B2 VSS 6 3 1 4
c1 1 VSS 0.00749589f
c2 3 VSS 0.0465533f
c3 4 VSS 0.00488644f
r1 7 8 5.88804 $w=1.3e-08 $l=2.53e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1097 $X2=0.1890 $Y2=0.1350
r2 6 7 3.90593 $w=1.3e-08 $l=1.67e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0930 $X2=0.1890 $Y2=0.1097
r3 6 4 2.73998 $w=1.3e-08 $l=1.18e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0930 $X2=0.1890 $Y2=0.0812
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AO222x2_ASAP7_75t_R%A1 VSS 8 3 1 4
c1 1 VSS 0.00748825f
c2 3 VSS 0.0463903f
c3 4 VSS 0.0057318f
r1 8 7 0.408082 $w=1.3e-08 $l=1.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1470 $X2=0.4050 $Y2=0.1452
r2 6 7 2.39019 $w=1.3e-08 $l=1.02e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1452
r3 4 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0980 $X2=0.4050 $Y2=0.1350
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r5 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
.ends

.subckt PM_AO222x2_ASAP7_75t_R%NET17 VSS 16 17 31 33 10 1 11 2 12 3 13
c1 1 VSS 0.0051357f
c2 2 VSS 0.00458232f
c3 3 VSS 0.00566825f
c4 10 VSS 0.00223963f
c5 11 VSS 0.00219195f
c6 12 VSS 0.00312799f
c7 13 VSS 0.0212428f
r1 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2680 $Y2=0.2025
r2 33 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r3 31 30 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r4 10 30 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r5 3 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.2340
r6 1 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r7 27 28 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2315
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r8 26 27 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2000
+ $Y=0.2340 $X2=0.2315 $Y2=0.2340
r9 25 26 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.2000 $Y2=0.2340
r10 23 24 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2340 $X2=0.0925 $Y2=0.2340
r11 21 24 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1240
+ $Y=0.2340 $X2=0.0925 $Y2=0.2340
r12 20 21 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1240 $Y2=0.2340
r13 19 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1755
+ $Y=0.2340 $X2=0.1890 $Y2=0.2340
r14 18 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r15 13 18 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r16 13 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r17 2 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r18 16 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r19 2 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r20 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r21 17 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r22 1 10 1e-05
.ends

.subckt PM_AO222x2_ASAP7_75t_R%A2 VSS 6 3 4 1
c1 1 VSS 0.00770744f
c2 3 VSS 0.0835176f
c3 4 VSS 0.0057813f
r1 7 8 6.47102 $w=1.3e-08 $l=2.78e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1072 $X2=0.4590 $Y2=0.1350
r2 6 7 4.4889 $w=1.3e-08 $l=1.92e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0880 $X2=0.4590 $Y2=0.1072
r3 6 4 2.15701 $w=1.3e-08 $l=9.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0880 $X2=0.4590 $Y2=0.0787
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1350
+ $X2=0.4590 $Y2=0.1350
.ends

.subckt PM_AO222x2_ASAP7_75t_R%NET18 VSS 16 17 31 32 7 1 9 8 11 2
c1 1 VSS 0.00327391f
c2 2 VSS 0.00989667f
c3 7 VSS 0.00248245f
c4 8 VSS 0.00484865f
c5 9 VSS 0.00313808f
c6 10 VSS 0.000841271f
c7 11 VSS 0.0116697f
c8 12 VSS 0.00092227f
c9 13 VSS 0.00294733f
r1 32 30 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r2 2 30 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r4 31 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r5 2 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.2340
r6 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4185
+ $Y=0.2340 $X2=0.4320 $Y2=0.2340
r7 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.2340 $X2=0.4185 $Y2=0.2340
r8 11 13 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3780 $Y=0.2340 $X2=0.3510 $Y2=0.2340
r9 11 24 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.4050 $Y2=0.2340
r10 10 23 2.45586 $w=1.44e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.2160 $X2=0.3510 $Y2=0.2035
r11 10 13 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.2160 $X2=0.3510 $Y2=0.2340
r12 12 23 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1945 $X2=0.3510 $Y2=0.2035
r13 22 23 7.11966 $w=1.35385e-08 $l=3.8396e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3130 $Y=0.1980 $X2=0.3510 $Y2=0.2035
r14 21 22 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2680
+ $Y=0.1980 $X2=0.3130 $Y2=0.1980
r15 20 21 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1980 $X2=0.2680 $Y2=0.1980
r16 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.1980 $X2=0.2430 $Y2=0.1980
r17 18 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1980 $X2=0.2295 $Y2=0.1980
r18 9 18 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2045
+ $Y=0.1980 $X2=0.2160 $Y2=0.1980
r19 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.1980
r20 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r21 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r22 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r23 16 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
.ends


*
.SUBCKT AO222x2_ASAP7_75t_R VSS VDD C1 C2 B2 B1 A1 A2 Y
*
* VSS VSS
* VDD VDD
* C1 C1
* C2 C2
* B2 B2
* B1 B1
* A1 A1
* A2 A2
* Y Y
*
*

MM10 N_MM10_d N_MM10_g N_MM10_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 N_MM11_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM14 N_MM14_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM13 N_MM13_d N_MM1_g N_MM13_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM0_g N_MM6_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM8_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9@2 N_MM9@2_d N_MM8@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM10_g N_MM2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM11_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g N_MM4_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM8_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8@2 N_MM8@2_d N_MM8@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AO222x2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AO222x2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AO222x2_ASAP7_75t_R%NET36 VSS N_MM10_s N_MM11_d N_NET36_1
+ PM_AO222x2_ASAP7_75t_R%NET36
cc_1 N_NET36_1 N_MM10_g 0.0173484f
cc_2 N_NET36_1 N_MM11_g 0.0174365f
x_PM_AO222x2_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_AO222x2_ASAP7_75t_R%noxref_21
cc_3 N_noxref_21_1 N_MM0_g 0.00140287f
cc_4 N_noxref_21_1 N_noxref_19_1 0.00767306f
cc_5 N_noxref_21_1 N_noxref_20_1 0.00123597f
x_PM_AO222x2_ASAP7_75t_R%NET37 VSS N_MM14_d N_MM13_s N_NET37_1
+ PM_AO222x2_ASAP7_75t_R%NET37
cc_6 N_NET37_1 N_MM4_g 0.0172226f
cc_7 N_NET37_1 N_MM1_g 0.0173091f
x_PM_AO222x2_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_AO222x2_ASAP7_75t_R%noxref_19
cc_8 N_noxref_19_1 N_MM1_g 0.0013908f
cc_9 N_noxref_19_1 N_NET17_12 0.0357683f
cc_10 N_noxref_19_1 N_noxref_18_1 0.00123731f
x_PM_AO222x2_ASAP7_75t_R%NET38 VSS N_MM6_s N_MM7_d N_NET38_1
+ PM_AO222x2_ASAP7_75t_R%NET38
cc_11 N_NET38_1 N_MM0_g 0.0172413f
cc_12 N_NET38_1 N_MM3_g 0.0172902f
x_PM_AO222x2_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_AO222x2_ASAP7_75t_R%noxref_23
cc_13 N_noxref_23_1 N_MM8@2_g 0.00147486f
cc_14 N_noxref_23_1 N_Y_8 0.000840977f
cc_15 N_noxref_23_1 N_noxref_22_1 0.00177678f
x_PM_AO222x2_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_AO222x2_ASAP7_75t_R%noxref_16
cc_16 N_noxref_16_1 N_MM10_g 0.00146754f
cc_17 N_noxref_16_1 N_NET23_21 0.000330984f
cc_18 N_noxref_16_1 N_NET23_3 0.000501075f
cc_19 N_noxref_16_1 N_NET23_17 0.0372086f
cc_20 N_noxref_16_1 N_NET17_10 0.000465692f
x_PM_AO222x2_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_AO222x2_ASAP7_75t_R%noxref_22
cc_21 N_noxref_22_1 N_MM8@2_g 0.00146748f
cc_22 N_noxref_22_1 N_Y_7 0.000842356f
x_PM_AO222x2_ASAP7_75t_R%Y VSS Y N_MM9_d N_MM9@2_d N_MM8_d N_MM8@2_d N_Y_7
+ N_Y_8 N_Y_12 N_Y_13 N_Y_10 N_Y_2 N_Y_1 PM_AO222x2_ASAP7_75t_R%Y
cc_23 N_Y_7 N_NET23_28 0.000179643f
cc_24 N_Y_7 N_NET23_29 0.000233849f
cc_25 N_Y_7 N_NET23_25 0.000350396f
cc_26 N_Y_7 N_NET23_24 0.00053784f
cc_27 N_Y_7 N_NET23_1 0.000883012f
cc_28 N_Y_8 N_MM8@2_g 0.0310268f
cc_29 N_Y_12 N_NET23_25 0.00104186f
cc_30 N_Y_13 N_NET23_28 0.00119926f
cc_31 N_Y_10 N_NET23_25 0.00145434f
cc_32 N_Y_2 N_MM8@2_g 0.00213081f
cc_33 N_Y_1 N_MM8@2_g 0.00218872f
cc_34 N_Y_10 N_NET23_24 0.00296635f
cc_35 N_Y_8 N_NET23_1 0.00443089f
cc_36 N_Y_7 N_MM8_g 0.0372607f
cc_37 N_Y_7 N_MM8@2_g 0.0684158f
x_PM_AO222x2_ASAP7_75t_R%C2 VSS C2 N_MM11_g N_C2_1 N_C2_4
+ PM_AO222x2_ASAP7_75t_R%C2
cc_38 N_C2_1 N_C1_1 0.00119807f
cc_39 N_C2_4 N_C1_4 0.00340994f
cc_40 N_MM11_g N_MM10_g 0.00590171f
x_PM_AO222x2_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_AO222x2_ASAP7_75t_R%noxref_20
cc_41 N_noxref_20_1 N_MM0_g 0.00141681f
cc_42 N_noxref_20_1 N_NET23_6 0.000423609f
cc_43 N_noxref_20_1 N_NET23_19 0.0374222f
cc_44 N_noxref_20_1 N_noxref_18_1 0.00767799f
x_PM_AO222x2_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_AO222x2_ASAP7_75t_R%noxref_17
cc_45 N_noxref_17_1 N_MM10_g 0.00144878f
cc_46 N_noxref_17_1 N_NET23_21 0.000256364f
cc_47 N_noxref_17_1 N_NET23_20 0.00106305f
cc_48 N_noxref_17_1 N_NET17_10 0.0360908f
cc_49 N_noxref_17_1 N_noxref_16_1 0.00175581f
x_PM_AO222x2_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_AO222x2_ASAP7_75t_R%noxref_18
cc_50 N_noxref_18_1 N_MM1_g 0.0014197f
cc_51 N_noxref_18_1 N_NET23_5 0.0004247f
cc_52 N_noxref_18_1 N_NET23_18 0.0372223f
x_PM_AO222x2_ASAP7_75t_R%C1 VSS C1 N_MM10_g N_C1_1 N_C1_4
+ PM_AO222x2_ASAP7_75t_R%C1
x_PM_AO222x2_ASAP7_75t_R%NET23 VSS N_MM8_g N_MM8@2_g N_MM6_d N_MM13_d N_MM10_d
+ N_MM2_d N_MM5_d N_NET23_20 N_NET23_3 N_NET23_4 N_NET23_23 N_NET23_22
+ N_NET23_21 N_NET23_17 N_NET23_18 N_NET23_5 N_NET23_6 N_NET23_19 N_NET23_25
+ N_NET23_1 N_NET23_24 N_NET23_29 N_NET23_27 N_NET23_28
+ PM_AO222x2_ASAP7_75t_R%NET23
cc_53 N_NET23_20 N_MM10_g 0.0157087f
cc_54 N_NET23_3 N_C1_1 0.000899013f
cc_55 N_NET23_4 N_MM10_g 0.000926567f
cc_56 N_NET23_23 N_C1_4 0.00121387f
cc_57 N_NET23_22 N_C1_4 0.00123453f
cc_58 N_NET23_3 N_MM10_g 0.0017316f
cc_59 N_NET23_20 N_C1_1 0.00181591f
cc_60 N_NET23_21 N_C1_4 0.00594737f
cc_61 N_NET23_17 N_MM10_g 0.0547443f
cc_62 N_NET23_3 N_MM11_g 0.000244211f
cc_63 N_NET23_4 N_MM11_g 0.00127355f
cc_64 N_NET23_23 N_C2_4 0.00061122f
cc_65 N_NET23_20 N_C2_1 0.000852233f
cc_66 N_NET23_22 N_C2_4 0.00130936f
cc_67 N_NET23_4 N_C2_4 0.00213719f
cc_68 N_NET23_20 N_MM11_g 0.0353362f
cc_69 N_NET23_18 N_B2_4 0.00039697f
cc_70 N_NET23_5 N_B2_4 0.000246638f
cc_71 N_NET23_22 N_B2_4 0.00317495f
cc_72 N_NET23_5 N_MM1_g 0.0021851f
cc_73 N_NET23_18 N_B1_1 0.000936366f
cc_74 N_NET23_22 N_B1_4 0.00156424f
cc_75 N_NET23_5 N_B1_4 0.00234494f
cc_76 N_NET23_18 N_MM1_g 0.0357418f
cc_77 N_NET23_6 N_MM0_g 0.00235936f
cc_78 N_NET23_19 N_A1_1 0.000919563f
cc_79 N_NET23_22 N_A1_4 0.001567f
cc_80 N_NET23_6 N_A1_4 0.00249379f
cc_81 N_NET23_19 N_MM0_g 0.0358921f
cc_82 N_NET23_6 N_A2_4 0.000246854f
cc_83 N_NET23_25 N_A2_4 0.000336179f
cc_84 N_NET23_22 N_A2_4 0.00101751f
cc_85 N_NET23_1 N_A2_1 0.0010349f
cc_86 N_NET23_24 N_A2_4 0.00243435f
cc_87 N_MM8_g N_MM3_g 0.0035709f
cc_88 N_NET23_29 N_A2_4 0.00666672f
x_PM_AO222x2_ASAP7_75t_R%B1 VSS B1 N_MM1_g N_B1_1 N_B1_4
+ PM_AO222x2_ASAP7_75t_R%B1
cc_89 N_B1_1 N_B2_1 0.00117036f
cc_90 N_B1_4 N_B2_4 0.0033888f
cc_91 N_MM1_g N_MM4_g 0.00581359f
x_PM_AO222x2_ASAP7_75t_R%B2 VSS B2 N_MM4_g N_B2_1 N_B2_4
+ PM_AO222x2_ASAP7_75t_R%B2
cc_92 N_B2_1 N_C2_4 0.000819873f
cc_93 N_MM4_g N_MM11_g 0.0032683f
cc_94 N_B2_4 N_C2_4 0.00414156f
x_PM_AO222x2_ASAP7_75t_R%A1 VSS A1 N_MM0_g N_A1_1 N_A1_4
+ PM_AO222x2_ASAP7_75t_R%A1
x_PM_AO222x2_ASAP7_75t_R%NET17 VSS N_MM4_d N_MM5_s N_MM2_s N_MM1_d N_NET17_10
+ N_NET17_1 N_NET17_11 N_NET17_2 N_NET17_12 N_NET17_3 N_NET17_13
+ PM_AO222x2_ASAP7_75t_R%NET17
cc_95 N_NET17_10 N_C1_1 0.000747042f
cc_96 N_NET17_1 N_MM10_g 0.00104108f
cc_97 N_NET17_10 N_MM10_g 0.0343837f
cc_98 N_NET17_11 N_C2_1 0.000743588f
cc_99 N_NET17_2 N_MM11_g 0.000938037f
cc_100 N_NET17_11 N_MM11_g 0.0344888f
cc_101 N_NET17_11 N_B2_1 0.00073232f
cc_102 N_NET17_2 N_MM4_g 0.000939978f
cc_103 N_NET17_11 N_MM4_g 0.0345938f
cc_104 N_NET17_12 N_B1_1 0.000725454f
cc_105 N_NET17_3 N_MM1_g 0.00108737f
cc_106 N_NET17_12 N_MM1_g 0.0344267f
cc_107 N_NET17_13 N_NET23_17 9.63893e-20
cc_108 N_NET17_13 N_NET23_20 0.000100798f
cc_109 N_NET17_13 N_NET23_3 0.000136667f
cc_110 N_NET17_13 N_NET23_5 0.000146889f
cc_111 N_NET17_13 N_NET23_18 0.000421977f
cc_112 N_NET17_13 N_NET23_4 0.00121857f
cc_113 N_NET17_13 N_NET23_27 0.000446855f
cc_114 N_NET17_1 N_NET23_23 0.000555094f
cc_115 N_NET17_11 N_NET23_20 0.0016915f
cc_116 N_NET17_1 N_NET23_21 0.000638148f
cc_117 N_NET17_10 N_NET23_20 0.000779666f
cc_118 N_NET17_1 N_NET23_4 0.00249699f
cc_119 N_NET17_2 N_NET23_4 0.00416607f
cc_120 N_NET17_13 N_NET23_23 0.00889546f
x_PM_AO222x2_ASAP7_75t_R%A2 VSS A2 N_MM3_g N_A2_4 N_A2_1
+ PM_AO222x2_ASAP7_75t_R%A2
cc_121 N_MM3_g N_A1_1 0.00128876f
cc_122 N_A2_4 N_A1_4 0.00482619f
cc_123 N_MM3_g N_MM0_g 0.00585197f
x_PM_AO222x2_ASAP7_75t_R%NET18 VSS N_MM4_s N_MM1_s N_MM0_d N_MM3_d N_NET18_7
+ N_NET18_1 N_NET18_9 N_NET18_8 N_NET18_11 N_NET18_2
+ PM_AO222x2_ASAP7_75t_R%NET18
cc_124 N_NET18_7 N_B2_4 0.000615414f
cc_125 N_NET18_7 N_B2_1 0.0007582f
cc_126 N_NET18_1 N_B2_4 0.000789819f
cc_127 N_NET18_1 N_MM4_g 0.000870278f
cc_128 N_NET18_7 N_MM4_g 0.0337943f
cc_129 N_NET18_7 N_B1_1 0.000703257f
cc_130 N_NET18_1 N_MM1_g 0.000873721f
cc_131 N_NET18_9 N_B1_4 0.0014395f
cc_132 N_NET18_1 N_B1_4 0.0014797f
cc_133 N_NET18_7 N_MM1_g 0.0339846f
cc_134 N_NET18_8 N_A1_4 0.000519729f
cc_135 N_NET18_8 N_A1_1 0.000685043f
cc_136 N_NET18_11 N_A1_4 0.00108375f
cc_137 N_NET18_2 N_MM0_g 0.00117401f
cc_138 N_NET18_2 N_A1_4 0.0023874f
cc_139 N_NET18_8 N_MM0_g 0.034293f
cc_140 N_NET18_11 N_A2_4 0.000875629f
cc_141 N_NET18_2 N_MM3_g 0.00119138f
cc_142 N_NET18_2 N_A2_4 0.00151759f
cc_143 N_NET18_8 N_MM3_g 0.0345731f
cc_144 N_NET18_9 N_NET17_12 0.00062999f
cc_145 N_NET18_9 N_NET17_3 0.000715454f
cc_146 N_NET18_1 N_NET17_13 0.000773541f
cc_147 N_NET18_7 N_NET17_12 0.00112244f
cc_148 N_NET18_1 N_NET17_2 0.00133324f
cc_149 N_NET18_1 N_NET17_3 0.00499625f
cc_150 N_NET18_9 N_NET17_13 0.0103094f
*END of AO222x2_ASAP7_75t_R.pxi
.ENDS
** Design:	AO22x1_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AO22x1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AO22x1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AO22x1_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.0319521f
.ends

.subckt PM_AO22x1_ASAP7_75t_R%NET30 VSS 2 3 1
c1 1 VSS 0.000852956f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0540 $X2=0.1080 $Y2=0.0540
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0540 $X2=0.1080 $Y2=0.0540
.ends

.subckt PM_AO22x1_ASAP7_75t_R%NET29 VSS 2 3 1
c1 1 VSS 0.00086332f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0540 $X2=0.2160 $Y2=0.0540
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0540 $X2=0.2160 $Y2=0.0540
.ends

.subckt PM_AO22x1_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00497f
.ends

.subckt PM_AO22x1_ASAP7_75t_R%A1 VSS 16 3 6 1 5 9
c1 1 VSS 0.00185593f
c2 3 VSS 0.060793f
c3 4 VSS 0.00605364f
c4 5 VSS 0.00261393f
c5 6 VSS 0.00229654f
c6 7 VSS 0.00780057f
c7 8 VSS 0.00129726f
c8 9 VSS 0.00258984f
r1 9 17 5.29071 $w=1.46216e-08 $l=2.78e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1980 $X2=0.0270 $Y2=0.1702
r2 7 15 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0360 $X2=0.0270 $Y2=0.0540
r3 16 17 4.4889 $w=1.3e-08 $l=1.92e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1510 $X2=0.0270 $Y2=0.1702
r4 16 5 0.874462 $w=1.3e-08 $l=3.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1510 $X2=0.0270 $Y2=0.1472
r5 5 8 1.67627 $w=1.66735e-08 $l=1.22e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1472 $X2=0.0270 $Y2=0.1350
r6 14 15 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0720 $X2=0.0270 $Y2=0.0540
r7 4 8 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1035 $X2=0.0270 $Y2=0.1350
r8 4 14 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1035 $X2=0.0270 $Y2=0.0720
r9 8 13 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1350 $X2=0.0455 $Y2=0.1350
r10 6 11 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.0635
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r11 6 13 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0635
+ $Y=0.1350 $X2=0.0455 $Y2=0.1350
r12 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r13 1 11 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AO22x1_ASAP7_75t_R%B2 VSS 6 3 1 4
c1 1 VSS 0.00472714f
c2 3 VSS 0.00782837f
c3 4 VSS 0.00313039f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1207 $X2=0.1890 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1150 $X2=0.1890 $Y2=0.1207
r3 6 4 4.02252 $w=1.3e-08 $l=1.73e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1150 $X2=0.1890 $Y2=0.0977
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AO22x1_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.0421508f
.ends

.subckt PM_AO22x1_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.0421586f
.ends

.subckt PM_AO22x1_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.0317431f
.ends

.subckt PM_AO22x1_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.0048315f
.ends

.subckt PM_AO22x1_ASAP7_75t_R%B1 VSS 4 3 1 5
c1 1 VSS 0.00385095f
c2 3 VSS 0.034717f
c3 4 VSS 0.00272368f
c4 5 VSS 0.00335767f
r1 5 10 0.484711 $w=1.8e-08 $l=4.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.2382
+ $Y=0.0720 $X2=0.2430 $Y2=0.0720
r2 7 8 7.28718 $w=1.3e-08 $l=3.13e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1037 $X2=0.2430 $Y2=0.1350
r3 4 7 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0812 $X2=0.2430 $Y2=0.1037
r4 4 10 0.10932 $w=1.63333e-08 $l=9.2e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0812 $X2=0.2430 $Y2=0.0720
r5 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r6 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AO22x1_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00514326f
.ends

.subckt PM_AO22x1_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.00459526f
.ends

.subckt PM_AO22x1_ASAP7_75t_R%Y VSS 19 13 28 7 11 2 1 9 8
c1 1 VSS 0.00855657f
c2 2 VSS 0.00831471f
c3 7 VSS 0.00374334f
c4 8 VSS 0.00374139f
c5 9 VSS 0.00384723f
c6 10 VSS 0.00664546f
c7 11 VSS 0.00617973f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4300 $Y2=0.2025
r2 28 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r3 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.2340
r4 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4455 $Y2=0.2340
r5 11 22 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4590 $Y2=0.2160
r6 11 25 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.2340 $X2=0.4455 $Y2=0.2340
r7 21 22 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1755 $X2=0.4590 $Y2=0.2160
r8 20 21 7.98675 $w=1.3e-08 $l=3.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1412 $X2=0.4590 $Y2=0.1755
r9 19 20 0.757867 $w=1.3e-08 $l=3.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1380 $X2=0.4590 $Y2=0.1412
r10 19 18 1.45744 $w=1.3e-08 $l=6.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1380 $X2=0.4590 $Y2=0.1317
r11 9 17 10.3626 $w=1.39091e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0855 $X2=0.4590 $Y2=0.0360
r12 9 18 10.785 $w=1.3e-08 $l=4.62e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0855 $X2=0.4590 $Y2=0.1317
r13 16 17 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4455 $Y=0.0360 $X2=0.4590 $Y2=0.0360
r14 15 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4455 $Y2=0.0360
r15 14 15 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4210
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r16 10 14 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4185
+ $Y=0.0360 $X2=0.4210 $Y2=0.0360
r17 1 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4320 $Y2=0.0360
r18 7 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0675 $X2=0.4300 $Y2=0.0675
r19 13 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4175 $Y2=0.0675
.ends

.subckt PM_AO22x1_ASAP7_75t_R%A2 VSS 11 3 6 5 1 4
c1 1 VSS 0.00301978f
c2 3 VSS 0.0338922f
c3 4 VSS 0.00235886f
c4 5 VSS 0.00214524f
c5 6 VSS 0.00222748f
r1 6 12 1.20989 $w=1.73902e-08 $l=1.03e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1980 $X2=0.1350 $Y2=0.1877
r2 5 8 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.0720 $X2=0.1350 $Y2=0.1035
r3 11 12 0.408082 $w=1.3e-08 $l=1.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1860 $X2=0.1350 $Y2=0.1877
r4 11 10 2.62338 $w=1.3e-08 $l=1.13e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1860 $X2=0.1350 $Y2=0.1747
r5 9 10 4.83869 $w=1.3e-08 $l=2.07e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1540 $X2=0.1350 $Y2=0.1747
r6 4 8 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1035
r7 4 9 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1540
r8 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r9 1 4 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AO22x1_ASAP7_75t_R%NET13 VSS 15 31 32 34 1 13 10 11 2 3 12
c1 1 VSS 0.00744776f
c2 2 VSS 0.00638366f
c3 3 VSS 0.00556441f
c4 10 VSS 0.00325146f
c5 11 VSS 0.00294458f
c6 12 VSS 0.00268101f
c7 13 VSS 0.0216511f
r1 12 3 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2160 $X2=0.2680 $Y2=0.2160
r2 34 12 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2160 $X2=0.2555 $Y2=0.2160
r3 32 30 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2160 $X2=0.1765 $Y2=0.2160
r4 2 30 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2160 $X2=0.1765 $Y2=0.2160
r5 11 2 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1620 $Y2=0.2160
r6 31 11 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r7 3 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2160
+ $X2=0.2700 $Y2=0.2340
r8 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r9 26 27 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2315
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r10 25 26 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2000
+ $Y=0.2340 $X2=0.2315 $Y2=0.2340
r11 24 25 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.2000 $Y2=0.2340
r12 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1755
+ $Y=0.2340 $X2=0.1890 $Y2=0.2340
r13 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r14 21 22 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r15 20 21 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.1255
+ $Y=0.2340 $X2=0.1485 $Y2=0.2340
r16 19 20 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1010
+ $Y=0.2340 $X2=0.1255 $Y2=0.2340
r17 18 19 5.13017 $w=1.3e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0790
+ $Y=0.2340 $X2=0.1010 $Y2=0.2340
r18 17 18 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0590
+ $Y=0.2340 $X2=0.0790 $Y2=0.2340
r19 16 17 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0500
+ $Y=0.2340 $X2=0.0590 $Y2=0.2340
r20 13 16 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.2340 $X2=0.0500 $Y2=0.2340
r21 1 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0500 $Y2=0.2340
r22 15 14 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r23 10 14 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r24 1 10 1e-05
.ends

.subckt PM_AO22x1_ASAP7_75t_R%NET18 VSS 9 43 44 47 48 13 3 12 10 11 4 14 17 19
+ 1 16
c1 1 VSS 0.00418041f
c2 3 VSS 0.00556338f
c3 4 VSS 0.00295305f
c4 9 VSS 0.0803318f
c5 10 VSS 0.00404978f
c6 11 VSS 0.00305203f
c7 12 VSS 0.0248172f
c8 13 VSS 0.00347889f
c9 14 VSS 0.00384268f
c10 15 VSS 0.00175743f
c11 16 VSS 0.00180214f
c12 17 VSS 0.00394544f
c13 18 VSS 0.000344393f
c14 19 VSS 0.00185729f
r1 48 46 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2160 $X2=0.2305 $Y2=0.2160
r2 4 46 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2160 $X2=0.2305 $Y2=0.2160
r3 11 4 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2160 $X2=0.2160 $Y2=0.2160
r4 47 11 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2160 $X2=0.2015 $Y2=0.2160
r5 44 42 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0540 $X2=0.1765 $Y2=0.0540
r6 3 42 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.0540 $X2=0.1765 $Y2=0.0540
r7 10 3 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1620 $Y2=0.0540
r8 43 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r9 4 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2160
+ $X2=0.2160 $Y2=0.1980
r10 3 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r11 39 40 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1980 $X2=0.2295 $Y2=0.1980
r12 37 40 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1980 $X2=0.2295 $Y2=0.1980
r13 36 37 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2680
+ $Y=0.1980 $X2=0.2430 $Y2=0.1980
r14 35 36 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.2855
+ $Y=0.1980 $X2=0.2680 $Y2=0.1980
r15 13 19 6.86231 $w=1.42329e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3145 $Y=0.1980 $X2=0.3510 $Y2=0.1980
r16 13 35 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.3145
+ $Y=0.1980 $X2=0.2855 $Y2=0.1980
r17 32 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r18 30 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r19 29 30 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2000
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r20 28 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2180
+ $Y=0.0360 $X2=0.2000 $Y2=0.0360
r21 27 28 9.91056 $w=1.3e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2605
+ $Y=0.0360 $X2=0.2180 $Y2=0.0360
r22 12 17 6.86231 $w=1.42329e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3145 $Y=0.0360 $X2=0.3510 $Y2=0.0360
r23 12 27 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3145
+ $Y=0.0360 $X2=0.2605 $Y2=0.0360
r24 19 26 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.1980 $X2=0.3510 $Y2=0.1765
r25 17 25 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0360 $X2=0.3510 $Y2=0.0540
r26 15 18 3.2503 $w=1.53684e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.1540 $X2=0.3510 $Y2=0.1350
r27 15 26 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1540 $X2=0.3510 $Y2=0.1765
r28 24 25 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0720 $X2=0.3510 $Y2=0.0540
r29 14 18 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.1035 $X2=0.3510 $Y2=0.1350
r30 14 24 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1035 $X2=0.3510 $Y2=0.0720
r31 16 21 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r32 16 18 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3780 $Y=0.1350 $X2=0.3510 $Y2=0.1350
r33 9 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r34 1 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
.ends


*
.SUBCKT AO22x1_ASAP7_75t_R VSS VDD A1 A2 B2 B1 Y
*
* VSS VSS
* VDD VDD
* A1 A1
* A2 A2
* B2 B2
* B1 B1
* Y Y
*
*

MM8 N_MM8_d N_MM8_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM6 N_MM6_d N_MM6_g N_MM6_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM7 N_MM7_d N_MM7_g N_MM7_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM9 N_MM9_d N_MM9_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM0 N_MM0_d N_MM0_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM8_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM6_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM7_g N_MM5_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM4 N_MM4_d N_MM9_g N_MM4_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1 N_MM1_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AO22x1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AO22x1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AO22x1_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_AO22x1_ASAP7_75t_R%noxref_12
cc_1 N_noxref_12_1 N_MM8_g 0.00460248f
x_PM_AO22x1_ASAP7_75t_R%NET30 VSS N_MM8_d N_MM6_s N_NET30_1
+ PM_AO22x1_ASAP7_75t_R%NET30
cc_2 N_NET30_1 N_MM8_g 0.0125072f
cc_3 N_NET30_1 N_MM6_g 0.0125729f
x_PM_AO22x1_ASAP7_75t_R%NET29 VSS N_MM7_s N_MM9_d N_NET29_1
+ PM_AO22x1_ASAP7_75t_R%NET29
cc_4 N_NET29_1 N_MM7_g 0.0125919f
cc_5 N_NET29_1 N_MM9_g 0.0127286f
x_PM_AO22x1_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_AO22x1_ASAP7_75t_R%noxref_13
cc_6 N_noxref_13_1 N_MM8_g 0.0044923f
cc_7 N_noxref_13_1 N_NET13_10 0.0270375f
cc_8 N_noxref_13_1 N_noxref_12_1 0.00205502f
x_PM_AO22x1_ASAP7_75t_R%A1 VSS A1 N_MM8_g N_A1_6 N_A1_1 N_A1_5 N_A1_9
+ PM_AO22x1_ASAP7_75t_R%A1
x_PM_AO22x1_ASAP7_75t_R%B2 VSS B2 N_MM7_g N_B2_1 N_B2_4 PM_AO22x1_ASAP7_75t_R%B2
cc_9 N_B2_1 N_MM6_g 0.000961944f
cc_10 N_B2_1 N_A2_1 0.0016438f
cc_11 N_B2_4 N_A2_4 0.00367387f
cc_12 N_MM7_g N_MM6_g 0.00798251f
x_PM_AO22x1_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_AO22x1_ASAP7_75t_R%noxref_16
cc_13 N_noxref_16_1 N_MM0_g 0.00175424f
cc_14 N_noxref_16_1 N_noxref_14_1 0.00771715f
cc_15 N_noxref_16_1 N_noxref_15_1 0.000471599f
x_PM_AO22x1_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_AO22x1_ASAP7_75t_R%noxref_17
cc_16 N_noxref_17_1 N_MM0_g 0.00174219f
cc_17 N_noxref_17_1 N_noxref_14_1 0.000472615f
cc_18 N_noxref_17_1 N_noxref_15_1 0.00769874f
cc_19 N_noxref_17_1 N_noxref_16_1 0.00123847f
x_PM_AO22x1_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_AO22x1_ASAP7_75t_R%noxref_14
cc_20 N_noxref_14_1 N_MM9_g 0.00368453f
cc_21 N_noxref_14_1 N_MM0_g 0.000534389f
x_PM_AO22x1_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_AO22x1_ASAP7_75t_R%noxref_18
cc_22 N_noxref_18_1 N_MM0_g 0.00145321f
cc_23 N_noxref_18_1 N_Y_7 0.0383747f
x_PM_AO22x1_ASAP7_75t_R%B1 VSS B1 N_MM9_g N_B1_1 N_B1_5 PM_AO22x1_ASAP7_75t_R%B1
cc_24 N_B1_1 N_MM7_g 0.000950699f
cc_25 N_B1_1 N_B2_1 0.00173244f
cc_26 N_B1 N_B2_4 0.00326866f
cc_27 N_MM9_g N_MM7_g 0.00915818f
x_PM_AO22x1_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_AO22x1_ASAP7_75t_R%noxref_15
cc_28 N_noxref_15_1 N_MM9_g 0.00360617f
cc_29 N_noxref_15_1 N_NET18_11 0.000634427f
cc_30 N_noxref_15_1 N_NET13_12 0.026626f
cc_31 N_noxref_15_1 N_noxref_14_1 0.00147317f
x_PM_AO22x1_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_AO22x1_ASAP7_75t_R%noxref_19
cc_32 N_noxref_19_1 N_MM0_g 0.00144894f
cc_33 N_noxref_19_1 N_Y_8 0.0385543f
cc_34 N_noxref_19_1 N_noxref_18_1 0.00177366f
x_PM_AO22x1_ASAP7_75t_R%Y VSS Y N_MM0_d N_MM1_d N_Y_7 N_Y_11 N_Y_2 N_Y_1 N_Y_9
+ N_Y_8 PM_AO22x1_ASAP7_75t_R%Y
cc_35 N_Y_7 N_NET18_14 0.000524446f
cc_36 N_Y_7 N_NET18_17 0.000546296f
cc_37 N_Y_11 N_NET18_19 0.000606888f
cc_38 N_Y_2 N_MM0_g 0.00117134f
cc_39 N_Y_1 N_MM0_g 0.00119169f
cc_40 N_Y_2 N_NET18_1 0.00121679f
cc_41 N_Y_7 N_NET18_1 0.00160378f
cc_42 N_Y_9 N_NET18_16 0.00374318f
cc_43 N_Y_8 N_MM0_g 0.0154557f
cc_44 N_Y_7 N_MM0_g 0.0550456f
x_PM_AO22x1_ASAP7_75t_R%A2 VSS A2 N_MM6_g N_A2_6 N_A2_5 N_A2_1 N_A2_4
+ PM_AO22x1_ASAP7_75t_R%A2
cc_45 N_A2_6 N_A1_6 0.000482767f
cc_46 N_A2_5 N_A1_6 0.0006329f
cc_47 N_A2_1 N_A1_1 0.0023585f
cc_48 N_A2_4 N_A1_6 0.00269042f
cc_49 N_MM6_g N_MM8_g 0.0101117f
x_PM_AO22x1_ASAP7_75t_R%NET13 VSS N_MM2_d N_MM3_d N_MM5_s N_MM4_s N_NET13_1
+ N_NET13_13 N_NET13_10 N_NET13_11 N_NET13_2 N_NET13_3 N_NET13_12
+ PM_AO22x1_ASAP7_75t_R%NET13
cc_50 N_NET13_1 N_A1_5 0.000386938f
cc_51 N_NET13_1 N_MM8_g 0.00119542f
cc_52 N_NET13_13 N_A1_9 0.00357482f
cc_53 N_NET13_10 N_MM8_g 0.0259582f
cc_54 N_NET13_11 N_A2_4 0.000544953f
cc_55 N_NET13_2 N_MM6_g 0.00072802f
cc_56 N_NET13_13 N_A2_6 0.00485088f
cc_57 N_NET13_11 N_MM6_g 0.0252583f
cc_58 N_NET13_2 N_MM7_g 0.000529911f
cc_59 N_NET13_11 N_MM7_g 0.0255434f
cc_60 N_NET13_3 N_MM9_g 0.000604788f
cc_61 N_NET13_12 N_MM9_g 0.025375f
cc_62 N_NET13_13 N_NET18_11 0.000924625f
cc_63 N_NET13_3 N_NET18_13 0.000599722f
cc_64 N_NET13_13 N_NET18_4 0.000743081f
cc_65 N_NET13_12 N_NET18_11 0.000837849f
cc_66 N_NET13_2 N_NET18_4 0.000975476f
cc_67 N_NET13_3 N_NET18_4 0.00380181f
cc_68 N_NET13_13 N_NET18_13 0.00973465f
x_PM_AO22x1_ASAP7_75t_R%NET18 VSS N_MM0_g N_MM6_d N_MM7_d N_MM5_d N_MM4_d
+ N_NET18_13 N_NET18_3 N_NET18_12 N_NET18_10 N_NET18_11 N_NET18_4 N_NET18_14
+ N_NET18_17 N_NET18_19 N_NET18_1 N_NET18_16 PM_AO22x1_ASAP7_75t_R%NET18
cc_69 N_NET18_13 N_MM6_g 0.000326882f
cc_70 N_NET18_3 N_A2_4 0.000648155f
cc_71 N_NET18_3 N_MM6_g 0.00103122f
cc_72 N_NET18_12 N_A2_5 0.0039845f
cc_73 N_NET18_10 N_MM6_g 0.026226f
cc_74 N_NET18_11 N_MM7_g 0.0112426f
cc_75 N_NET18_4 N_MM7_g 0.000410025f
cc_76 N_NET18_11 N_B2_1 0.000567908f
cc_77 N_NET18_13 N_B2_4 0.000587508f
cc_78 N_NET18_3 N_MM7_g 0.000948203f
cc_79 N_NET18_12 N_B2_4 0.00124156f
cc_80 N_NET18_3 N_B2_4 0.00231842f
cc_81 N_NET18_10 N_MM7_g 0.0398726f
cc_82 N_NET18_4 N_MM9_g 0.000725349f
cc_83 N_NET18_13 N_B1_1 0.000406645f
cc_84 N_NET18_11 N_B1_1 0.000547769f
cc_85 N_NET18_14 N_B1_5 0.000573118f
cc_86 N_NET18_13 N_B1 0.00360348f
cc_87 N_NET18_12 N_B1_5 0.00633237f
cc_88 N_NET18_11 N_MM9_g 0.0261181f
*END of AO22x1_ASAP7_75t_R.pxi
.ENDS
** Design:	AO22x2_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AO22x2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AO22x2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AO22x2_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.0430258f
.ends

.subckt PM_AO22x2_ASAP7_75t_R%NET29 VSS 2 3 1
c1 1 VSS 0.0010156f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2160 $Y2=0.0675
.ends

.subckt PM_AO22x2_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.0427357f
.ends

.subckt PM_AO22x2_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00714693f
.ends

.subckt PM_AO22x2_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.0423185f
.ends

.subckt PM_AO22x2_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.0423043f
.ends

.subckt PM_AO22x2_ASAP7_75t_R%Y VSS 22 16 17 31 32 7 8 11 2 1
c1 1 VSS 0.0104989f
c2 2 VSS 0.0104683f
c3 7 VSS 0.00455484f
c4 8 VSS 0.00454326f
c5 9 VSS 0.00972459f
c6 10 VSS 0.00976267f
c7 11 VSS 0.00758555f
c8 12 VSS 0.00348907f
c9 13 VSS 0.003492f
r1 32 30 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r2 2 30 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r4 31 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r5 2 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.2340
r6 26 27 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4725 $Y2=0.2340
r7 10 26 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4210
+ $Y=0.2340 $X2=0.4320 $Y2=0.2340
r8 13 25 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.2340 $X2=0.5130 $Y2=0.2160
r9 13 27 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.2340 $X2=0.4725 $Y2=0.2340
r10 24 25 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1755 $X2=0.5130 $Y2=0.2160
r11 23 24 7.98675 $w=1.3e-08 $l=3.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1412 $X2=0.5130 $Y2=0.1755
r12 22 23 0.757867 $w=1.3e-08 $l=3.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1380 $X2=0.5130 $Y2=0.1412
r13 22 21 1.45744 $w=1.3e-08 $l=6.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1380 $X2=0.5130 $Y2=0.1317
r14 11 12 9.89378 $w=1.47818e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.0855 $X2=0.5130 $Y2=0.0360
r15 11 21 10.785 $w=1.3e-08 $l=4.62e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0855 $X2=0.5130 $Y2=0.1317
r16 12 20 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.0360 $X2=0.4725 $Y2=0.0360
r17 19 20 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4725 $Y2=0.0360
r18 18 19 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4210
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r19 9 18 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4185
+ $Y=0.0360 $X2=0.4210 $Y2=0.0360
r20 1 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4320 $Y2=0.0360
r21 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r22 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r23 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0675 $X2=0.4320 $Y2=0.0675
r24 16 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4175 $Y2=0.0675
.ends

.subckt PM_AO22x2_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.0421789f
.ends

.subckt PM_AO22x2_ASAP7_75t_R%NET18 VSS 9 10 54 55 58 59 14 3 11 13 4 12 15 16
+ 1 17
c1 1 VSS 0.0091674f
c2 3 VSS 0.00630146f
c3 4 VSS 0.00300308f
c4 9 VSS 0.0814035f
c5 10 VSS 0.0807835f
c6 11 VSS 0.00578793f
c7 12 VSS 0.00487117f
c8 13 VSS 0.0259167f
c9 14 VSS 0.00425633f
c10 15 VSS 0.00447971f
c11 16 VSS 0.00210056f
c12 17 VSS 0.00275382f
c13 18 VSS 0.00370623f
c14 19 VSS 0.000465159f
c15 20 VSS 0.00191877f
r1 59 57 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r2 4 57 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r3 12 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r4 58 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r5 55 53 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r6 3 53 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r7 11 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r8 54 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1475 $Y2=0.0675
r9 4 50 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.1980
r10 3 43 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0675
+ $X2=0.1620 $Y2=0.0360
r11 50 51 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1980 $X2=0.2295 $Y2=0.1980
r12 48 51 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1980 $X2=0.2295 $Y2=0.1980
r13 47 48 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2680
+ $Y=0.1980 $X2=0.2430 $Y2=0.1980
r14 46 47 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.2855
+ $Y=0.1980 $X2=0.2680 $Y2=0.1980
r15 14 20 6.86231 $w=1.42329e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3145 $Y=0.1980 $X2=0.3510 $Y2=0.1980
r16 14 46 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.3145
+ $Y=0.1980 $X2=0.2855 $Y2=0.1980
r17 43 44 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r18 41 44 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r19 40 41 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2000
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r20 39 40 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2180
+ $Y=0.0360 $X2=0.2000 $Y2=0.0360
r21 38 39 9.91056 $w=1.3e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2605
+ $Y=0.0360 $X2=0.2180 $Y2=0.0360
r22 13 18 6.86231 $w=1.42329e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3145 $Y=0.0360 $X2=0.3510 $Y2=0.0360
r23 13 38 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3145
+ $Y=0.0360 $X2=0.2605 $Y2=0.0360
r24 20 37 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.1980 $X2=0.3510 $Y2=0.1765
r25 18 36 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0360 $X2=0.3510 $Y2=0.0540
r26 16 19 3.2503 $w=1.53684e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.1540 $X2=0.3510 $Y2=0.1350
r27 16 37 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1540 $X2=0.3510 $Y2=0.1765
r28 35 36 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0720 $X2=0.3510 $Y2=0.0540
r29 15 19 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.1035 $X2=0.3510 $Y2=0.1350
r30 15 35 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1035 $X2=0.3510 $Y2=0.0720
r31 10 29 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r32 17 31 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r33 17 19 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3780 $Y=0.1350 $X2=0.3510 $Y2=0.1350
r34 27 29 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4465 $Y=0.1350 $X2=0.4590 $Y2=0.1350
r35 26 27 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4320 $Y=0.1350 $X2=0.4465 $Y2=0.1350
r36 25 26 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4175 $Y=0.1350 $X2=0.4320 $Y2=0.1350
r37 23 25 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.4145 $Y=0.1350 $X2=0.4175 $Y2=0.1350
r38 22 23 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4145 $Y2=0.1350
r39 22 31 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
r40 1 22 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.3955
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r41 1 24 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.3955
+ $Y=0.1350 $X2=0.3945 $Y2=0.1350
r42 9 22 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4050 $Y2=0.1350
r43 9 24 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.4050 $Y=0.1350 $X2=0.3945 $Y2=0.1350
r44 9 25 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4175 $Y2=0.1350
.ends

.subckt PM_AO22x2_ASAP7_75t_R%B2 VSS 6 3 1 4
c1 1 VSS 0.00674429f
c2 3 VSS 0.00880404f
c3 4 VSS 0.00422582f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1207 $X2=0.1890 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1150 $X2=0.1890 $Y2=0.1207
r3 6 4 4.02252 $w=1.3e-08 $l=1.73e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1150 $X2=0.1890 $Y2=0.0977
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AO22x2_ASAP7_75t_R%B1 VSS 4 3 1 5
c1 1 VSS 0.00679141f
c2 3 VSS 0.0461622f
c3 4 VSS 0.00391515f
c4 5 VSS 0.00445819f
r1 5 10 0.484711 $w=1.8e-08 $l=4.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.2382
+ $Y=0.0720 $X2=0.2430 $Y2=0.0720
r2 7 8 7.28718 $w=1.3e-08 $l=3.13e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1037 $X2=0.2430 $Y2=0.1350
r3 4 7 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0812 $X2=0.2430 $Y2=0.1037
r4 4 10 0.10932 $w=1.63333e-08 $l=9.2e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0812 $X2=0.2430 $Y2=0.0720
r5 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r6 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AO22x2_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00617749f
.ends

.subckt PM_AO22x2_ASAP7_75t_R%NET30 VSS 2 3 1
c1 1 VSS 0.0010141f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_AO22x2_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.0419296f
.ends

.subckt PM_AO22x2_ASAP7_75t_R%NET13 VSS 15 31 32 34 1 10 13 2 11 12 3
c1 1 VSS 0.00832609f
c2 2 VSS 0.00703848f
c3 3 VSS 0.00579203f
c4 10 VSS 0.00371425f
c5 11 VSS 0.00324472f
c6 12 VSS 0.00298228f
c7 13 VSS 0.0222674f
r1 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2680 $Y2=0.2025
r2 34 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r3 32 30 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r4 2 30 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r5 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r6 31 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r7 3 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.2340
r8 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r9 26 27 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2315
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r10 25 26 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2000
+ $Y=0.2340 $X2=0.2315 $Y2=0.2340
r11 24 25 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.2000 $Y2=0.2340
r12 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1755
+ $Y=0.2340 $X2=0.1890 $Y2=0.2340
r13 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r14 21 22 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r15 20 21 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.1255
+ $Y=0.2340 $X2=0.1485 $Y2=0.2340
r16 19 20 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1010
+ $Y=0.2340 $X2=0.1255 $Y2=0.2340
r17 18 19 5.13017 $w=1.3e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0790
+ $Y=0.2340 $X2=0.1010 $Y2=0.2340
r18 17 18 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0590
+ $Y=0.2340 $X2=0.0790 $Y2=0.2340
r19 16 17 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0500
+ $Y=0.2340 $X2=0.0590 $Y2=0.2340
r20 13 16 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.2340 $X2=0.0500 $Y2=0.2340
r21 1 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0500 $Y2=0.2340
r22 15 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r23 10 14 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r24 1 10 1e-05
.ends

.subckt PM_AO22x2_ASAP7_75t_R%A1 VSS 16 3 6 1 5 9
c1 1 VSS 0.0043779f
c2 3 VSS 0.082167f
c3 4 VSS 0.00738487f
c4 5 VSS 0.00307869f
c5 6 VSS 0.00262325f
c6 7 VSS 0.00840188f
c7 8 VSS 0.00155342f
c8 9 VSS 0.00290311f
r1 9 17 5.29071 $w=1.46216e-08 $l=2.78e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1980 $X2=0.0270 $Y2=0.1702
r2 7 15 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0360 $X2=0.0270 $Y2=0.0540
r3 16 17 4.4889 $w=1.3e-08 $l=1.92e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1510 $X2=0.0270 $Y2=0.1702
r4 16 5 0.874462 $w=1.3e-08 $l=3.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1510 $X2=0.0270 $Y2=0.1472
r5 5 8 1.67627 $w=1.66735e-08 $l=1.22e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1472 $X2=0.0270 $Y2=0.1350
r6 14 15 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0720 $X2=0.0270 $Y2=0.0540
r7 4 8 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1035 $X2=0.0270 $Y2=0.1350
r8 4 14 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1035 $X2=0.0270 $Y2=0.0720
r9 8 13 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1350 $X2=0.0455 $Y2=0.1350
r10 6 11 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.0635
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r11 6 13 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0635
+ $Y=0.1350 $X2=0.0455 $Y2=0.1350
r12 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r13 1 11 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AO22x2_ASAP7_75t_R%A2 VSS 11 3 5 1 4 6
c1 1 VSS 0.00536172f
c2 3 VSS 0.0451352f
c3 4 VSS 0.00330175f
c4 5 VSS 0.00290423f
c5 6 VSS 0.00301443f
r1 6 12 1.20989 $w=1.73902e-08 $l=1.03e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1980 $X2=0.1350 $Y2=0.1877
r2 5 8 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.0720 $X2=0.1350 $Y2=0.1035
r3 11 12 0.408082 $w=1.3e-08 $l=1.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1860 $X2=0.1350 $Y2=0.1877
r4 11 10 2.62338 $w=1.3e-08 $l=1.13e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1860 $X2=0.1350 $Y2=0.1747
r5 9 10 4.83869 $w=1.3e-08 $l=2.07e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1540 $X2=0.1350 $Y2=0.1747
r6 4 8 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1035
r7 4 9 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1540
r8 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r9 1 4 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends


*
.SUBCKT AO22x2_ASAP7_75t_R VSS VDD A1 A2 B2 B1 Y
*
* VSS VSS
* VDD VDD
* A1 A1
* A2 A2
* B2 B2
* B1 B1
* Y Y
*
*

MM8 N_MM8_d N_MM8_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM6_g N_MM6_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM7_g N_MM7_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM1_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@2 N_MM0@2_d N_MM1@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM8_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM6_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM7_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM9_g N_MM4_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1@2 N_MM1@2_d N_MM1@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AO22x2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AO22x2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AO22x2_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_AO22x2_ASAP7_75t_R%noxref_14
cc_1 N_noxref_14_1 N_MM9_g 0.00145657f
x_PM_AO22x2_ASAP7_75t_R%NET29 VSS N_MM7_s N_MM9_d N_NET29_1
+ PM_AO22x2_ASAP7_75t_R%NET29
cc_2 N_NET29_1 N_MM7_g 0.0172327f
cc_3 N_NET29_1 N_MM9_g 0.0173295f
x_PM_AO22x2_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_AO22x2_ASAP7_75t_R%noxref_16
cc_4 N_noxref_16_1 N_MM1_g 0.00177622f
cc_5 N_noxref_16_1 N_noxref_14_1 0.00765238f
x_PM_AO22x2_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_AO22x2_ASAP7_75t_R%noxref_15
cc_6 N_noxref_15_1 N_MM9_g 0.00139881f
cc_7 N_noxref_15_1 N_NET13_12 0.0359675f
cc_8 N_noxref_15_1 N_noxref_14_1 0.00124677f
x_PM_AO22x2_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_AO22x2_ASAP7_75t_R%noxref_18
cc_9 N_noxref_18_1 N_MM1@2_g 0.00146805f
cc_10 N_noxref_18_1 N_Y_7 0.000843573f
x_PM_AO22x2_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_AO22x2_ASAP7_75t_R%noxref_19
cc_11 N_noxref_19_1 N_MM1@2_g 0.00146658f
cc_12 N_noxref_19_1 N_Y_8 0.000836839f
cc_13 N_noxref_19_1 N_noxref_18_1 0.00177453f
x_PM_AO22x2_ASAP7_75t_R%Y VSS Y N_MM0_d N_MM0@2_d N_MM1_d N_MM1@2_d N_Y_7 N_Y_8
+ N_Y_11 N_Y_2 N_Y_1 PM_AO22x2_ASAP7_75t_R%Y
cc_14 N_Y_7 N_NET18_16 0.000245682f
cc_15 N_Y_7 N_NET18_15 0.000470922f
cc_16 N_Y_7 N_NET18_1 0.000645043f
cc_17 N_Y_8 N_MM1@2_g 0.030891f
cc_18 N_Y_11 N_NET18_1 0.000928226f
cc_19 N_Y_2 N_NET18_17 0.00109787f
cc_20 N_Y_1 N_MM1@2_g 0.00208413f
cc_21 N_Y_2 N_MM1@2_g 0.00212939f
cc_22 N_Y_8 N_NET18_1 0.00518076f
cc_23 N_Y_7 N_MM1_g 0.0372056f
cc_24 N_Y_7 N_MM1@2_g 0.0700875f
x_PM_AO22x2_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_AO22x2_ASAP7_75t_R%noxref_17
cc_25 N_noxref_17_1 N_MM1_g 0.00175501f
cc_26 N_noxref_17_1 N_NET13_12 0.00053554f
cc_27 N_noxref_17_1 N_noxref_15_1 0.00765898f
cc_28 N_noxref_17_1 N_noxref_16_1 0.00124037f
x_PM_AO22x2_ASAP7_75t_R%NET18 VSS N_MM1_g N_MM1@2_g N_MM6_d N_MM7_d N_MM5_d
+ N_MM4_d N_NET18_14 N_NET18_3 N_NET18_11 N_NET18_13 N_NET18_4 N_NET18_12
+ N_NET18_15 N_NET18_16 N_NET18_1 N_NET18_17 PM_AO22x2_ASAP7_75t_R%NET18
cc_29 N_NET18_14 N_MM6_g 0.000336581f
cc_30 N_NET18_3 N_A2_4 0.000820783f
cc_31 N_NET18_11 N_A2_1 0.000857627f
cc_32 N_NET18_3 N_MM6_g 0.00164761f
cc_33 N_NET18_13 N_A2_5 0.00415586f
cc_34 N_NET18_11 N_MM6_g 0.035885f
cc_35 N_NET18_4 N_B2_1 0.000528936f
cc_36 N_NET18_14 N_B2_4 0.000623368f
cc_37 N_NET18_4 N_MM7_g 0.000916962f
cc_38 N_NET18_13 N_B2_4 0.00118618f
cc_39 N_NET18_12 N_B2_1 0.00151043f
cc_40 N_NET18_3 N_MM7_g 0.00155074f
cc_41 N_NET18_3 N_B2_4 0.00261074f
cc_42 N_NET18_12 N_MM7_g 0.0150892f
cc_43 N_NET18_11 N_MM7_g 0.0550497f
cc_44 N_NET18_3 N_MM9_g 0.000242662f
cc_45 N_NET18_4 N_B1_1 0.000510677f
cc_46 N_NET18_15 N_B1_5 0.000514406f
cc_47 N_NET18_4 N_MM9_g 0.000927978f
cc_48 N_NET18_12 N_B1_1 0.00100797f
cc_49 N_NET18_14 N_B1 0.00355481f
cc_50 N_NET18_13 N_B1_5 0.00614373f
cc_51 N_NET18_12 N_MM9_g 0.0355864f
x_PM_AO22x2_ASAP7_75t_R%B2 VSS B2 N_MM7_g N_B2_1 N_B2_4 PM_AO22x2_ASAP7_75t_R%B2
cc_52 N_B2_1 N_A2_1 0.000849322f
cc_53 N_MM7_g N_MM6_g 0.00327732f
cc_54 N_B2_4 N_A2_4 0.00474689f
x_PM_AO22x2_ASAP7_75t_R%B1 VSS B1 N_MM9_g N_B1_1 N_B1_5 PM_AO22x2_ASAP7_75t_R%B1
cc_55 N_B1_1 N_B2_1 0.00126048f
cc_56 N_B1 N_B2_4 0.00325993f
cc_57 N_MM9_g N_MM7_g 0.00622359f
x_PM_AO22x2_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_AO22x2_ASAP7_75t_R%noxref_13
cc_58 N_noxref_13_1 N_MM8_g 0.00215013f
cc_59 N_noxref_13_1 N_NET13_10 0.0362956f
cc_60 N_noxref_13_1 N_noxref_12_1 0.00176447f
x_PM_AO22x2_ASAP7_75t_R%NET30 VSS N_MM8_d N_MM6_s N_NET30_1
+ PM_AO22x2_ASAP7_75t_R%NET30
cc_61 N_NET30_1 N_MM8_g 0.0171873f
cc_62 N_NET30_1 N_MM6_g 0.0172802f
x_PM_AO22x2_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_AO22x2_ASAP7_75t_R%noxref_12
cc_63 N_noxref_12_1 N_MM8_g 0.00224354f
cc_64 N_noxref_12_1 N_NET13_10 0.000478167f
x_PM_AO22x2_ASAP7_75t_R%NET13 VSS N_MM2_d N_MM3_d N_MM5_s N_MM4_s N_NET13_1
+ N_NET13_10 N_NET13_13 N_NET13_2 N_NET13_11 N_NET13_12 N_NET13_3
+ PM_AO22x2_ASAP7_75t_R%NET13
cc_65 N_NET13_1 N_A1_5 0.000537662f
cc_66 N_NET13_10 N_A1_1 0.000756499f
cc_67 N_NET13_1 N_MM8_g 0.00199235f
cc_68 N_NET13_13 N_A1_9 0.00360657f
cc_69 N_NET13_10 N_MM8_g 0.0353181f
cc_70 N_NET13_2 N_A2_4 0.000673429f
cc_71 N_NET13_2 N_MM6_g 0.00125962f
cc_72 N_NET13_13 N_A2_6 0.00474843f
cc_73 N_NET13_11 N_MM6_g 0.0348799f
cc_74 N_NET13_11 N_B2_1 0.000735104f
cc_75 N_NET13_2 N_MM7_g 0.000943013f
cc_76 N_NET13_11 N_MM7_g 0.0346702f
cc_77 N_NET13_12 N_B1_1 0.000910324f
cc_78 N_NET13_3 N_MM9_g 0.00109059f
cc_79 N_NET13_12 N_MM9_g 0.0346418f
cc_80 N_NET13_13 N_NET18_12 0.000599372f
cc_81 N_NET13_12 N_NET18_12 0.00179139f
cc_82 N_NET13_3 N_NET18_14 0.000768106f
cc_83 N_NET13_13 N_NET18_4 0.000771165f
cc_84 N_NET13_2 N_NET18_4 0.00137093f
cc_85 N_NET13_3 N_NET18_4 0.00508759f
cc_86 N_NET13_13 N_NET18_14 0.0103279f
x_PM_AO22x2_ASAP7_75t_R%A1 VSS A1 N_MM8_g N_A1_6 N_A1_1 N_A1_5 N_A1_9
+ PM_AO22x2_ASAP7_75t_R%A1
x_PM_AO22x2_ASAP7_75t_R%A2 VSS A2 N_MM6_g N_A2_5 N_A2_1 N_A2_4 N_A2_6
+ PM_AO22x2_ASAP7_75t_R%A2
cc_87 N_A2_5 N_A1_6 0.000590073f
cc_88 N_A2_1 N_A1_1 0.00185199f
cc_89 N_A2_4 N_A1_6 0.00266578f
cc_90 N_MM6_g N_MM8_g 0.00671315f
*END of AO22x2_ASAP7_75t_R.pxi
.ENDS
** Design:	AO31x2_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AO31x2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AO31x2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AO31x2_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00647997f
.ends

.subckt PM_AO31x2_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.0417379f
.ends

.subckt PM_AO31x2_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.0418689f
.ends

.subckt PM_AO31x2_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.0430869f
.ends

.subckt PM_AO31x2_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.0426822f
.ends

.subckt PM_AO31x2_ASAP7_75t_R%Y VSS 22 16 17 30 31 7 10 8 1 11 2
c1 1 VSS 0.0104634f
c2 2 VSS 0.010491f
c3 7 VSS 0.00453069f
c4 8 VSS 0.00454845f
c5 9 VSS 0.00965576f
c6 10 VSS 0.00957322f
c7 11 VSS 0.00723613f
c8 12 VSS 0.00349749f
c9 13 VSS 0.00351871f
r1 31 29 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.2025 $X2=0.7705 $Y2=0.2025
r2 2 29 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7560 $Y=0.2025 $X2=0.7705 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7415 $Y=0.2025 $X2=0.7560 $Y2=0.2025
r4 30 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.2025 $X2=0.7415 $Y2=0.2025
r5 2 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7560 $Y=0.2025
+ $X2=0.7560 $Y2=0.2340
r6 26 27 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.2340 $X2=0.7810 $Y2=0.2340
r7 9 13 4.06404 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8125 $Y=0.2340 $X2=0.8370 $Y2=0.2340
r8 9 27 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.8125
+ $Y=0.2340 $X2=0.7810 $Y2=0.2340
r9 13 24 9.89378 $w=1.47818e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8370 $Y=0.2340 $X2=0.8370 $Y2=0.1845
r10 23 24 10.9016 $w=1.3e-08 $l=4.68e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1377 $X2=0.8370 $Y2=0.1845
r11 22 23 1.57403 $w=1.3e-08 $l=6.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1310 $X2=0.8370 $Y2=0.1377
r12 22 21 0.641272 $w=1.3e-08 $l=2.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.1310 $X2=0.8370 $Y2=0.1282
r13 11 12 9.89378 $w=1.47818e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8370 $Y=0.0855 $X2=0.8370 $Y2=0.0360
r14 11 21 9.96886 $w=1.3e-08 $l=4.27e-08 $layer=M1 $thickness=3.6e-08 $X=0.8370
+ $Y=0.0855 $X2=0.8370 $Y2=0.1282
r15 12 20 4.06404 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8370 $Y=0.0360 $X2=0.8125 $Y2=0.0360
r16 19 20 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.7810
+ $Y=0.0360 $X2=0.8125 $Y2=0.0360
r17 18 19 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.0360 $X2=0.7810 $Y2=0.0360
r18 10 18 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.7445
+ $Y=0.0360 $X2=0.7560 $Y2=0.0360
r19 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7560 $Y=0.0675
+ $X2=0.7560 $Y2=0.0360
r20 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.0675 $X2=0.7705 $Y2=0.0675
r21 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7560 $Y=0.0675 $X2=0.7705 $Y2=0.0675
r22 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7415 $Y=0.0675 $X2=0.7560 $Y2=0.0675
r23 16 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.0675 $X2=0.7415 $Y2=0.0675
.ends

.subckt PM_AO31x2_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.0422995f
.ends

.subckt PM_AO31x2_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.0422996f
.ends

.subckt PM_AO31x2_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.00700425f
.ends

.subckt PM_AO31x2_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.00769391f
.ends

.subckt PM_AO31x2_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.0421185f
.ends

.subckt PM_AO31x2_ASAP7_75t_R%A1 VSS 21 3 4 9 1 7 6 8
c1 1 VSS 0.0100827f
c2 3 VSS 0.0456744f
c3 4 VSS 0.0459728f
c4 5 VSS 0.00347664f
c5 6 VSS 0.00327489f
c6 7 VSS 0.00399078f
c7 8 VSS 0.00327299f
c8 9 VSS 0.00390454f
r1 7 24 1.38478 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1620 $X2=0.5130 $Y2=0.1510
r2 5 8 4.18063 $w=1.6528e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1330 $X2=0.5130 $Y2=0.1080
r3 5 24 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1330 $X2=0.5130 $Y2=0.1510
r4 6 23 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5400 $Y=0.1080 $X2=0.5670 $Y2=0.1080
r5 6 8 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1080 $X2=0.5130 $Y2=0.1080
r6 21 9 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1215
r7 9 23 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.1215 $X2=0.5670 $Y2=0.1080
r8 4 17 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1350
r9 21 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1350
+ $X2=0.5670 $Y2=0.1350
r10 16 17 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.5575
+ $Y=0.1350 $X2=0.5670 $Y2=0.1350
r11 14 16 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.5545 $Y=0.1350 $X2=0.5575 $Y2=0.1350
r12 13 14 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5400 $Y=0.1350 $X2=0.5545 $Y2=0.1350
r13 12 13 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5255 $Y=0.1350 $X2=0.5400 $Y2=0.1350
r14 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r15 1 11 3.20232 $w=2.13909e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5020 $Y2=0.1350
r16 1 12 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5255 $Y2=0.1350
r17 3 11 0.905388 $w=2.07755e-07 $l=1.1e-08 $layer=LIG $thickness=5.52727e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5020 $Y2=0.1350
r18 3 12 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5255 $Y2=0.1350
.ends

.subckt PM_AO31x2_ASAP7_75t_R%A2 VSS 20 3 4 9 7 5 8 1 6
c1 1 VSS 0.0109653f
c2 3 VSS 0.0464065f
c3 4 VSS 0.0459171f
c4 5 VSS 0.00442319f
c5 6 VSS 0.00449276f
c6 7 VSS 0.00436193f
c7 8 VSS 0.00414479f
c8 9 VSS 0.00414635f
r1 8 28 1.38478 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1620 $X2=0.2970 $Y2=0.1510
r2 5 7 4.64944 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1330 $X2=0.2970 $Y2=0.1080
r3 5 28 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1330 $X2=0.2970 $Y2=0.1510
r4 7 25 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1080 $X2=0.3155 $Y2=0.1080
r5 24 25 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.3445
+ $Y=0.1080 $X2=0.3155 $Y2=0.1080
r6 6 22 4.64944 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3800
+ $Y=0.1080 $X2=0.4050 $Y2=0.1080
r7 6 24 8.27824 $w=1.3e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3800
+ $Y=0.1080 $X2=0.3445 $Y2=0.1080
r8 4 18 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r9 20 9 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1215
r10 9 22 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.1215 $X2=0.4050 $Y2=0.1080
r11 16 18 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4465 $Y=0.1350 $X2=0.4590 $Y2=0.1350
r12 15 16 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4320 $Y=0.1350 $X2=0.4465 $Y2=0.1350
r13 14 15 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4175 $Y=0.1350 $X2=0.4320 $Y2=0.1350
r14 12 14 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.4145 $Y=0.1350 $X2=0.4175 $Y2=0.1350
r15 11 12 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4145 $Y2=0.1350
r16 20 11 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
r17 1 11 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.3955
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r18 1 13 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.3955
+ $Y=0.1350 $X2=0.3945 $Y2=0.1350
r19 3 11 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4050 $Y2=0.1350
r20 3 13 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.4050 $Y=0.1350 $X2=0.3945 $Y2=0.1350
r21 3 14 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4175 $Y2=0.1350
.ends

.subckt PM_AO31x2_ASAP7_75t_R%NET30 VSS 15 33 34 36 2 1 13 11 10 3 12
c1 1 VSS 0.0038157f
c2 2 VSS 0.00318482f
c3 3 VSS 0.00395943f
c4 10 VSS 0.00289001f
c5 11 VSS 0.00215164f
c6 12 VSS 0.00291823f
c7 13 VSS 0.00274563f
r1 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.0675 $X2=0.5920 $Y2=0.0675
r2 36 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0675 $X2=0.5795 $Y2=0.0675
r3 34 32 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0675 $X2=0.5005 $Y2=0.0675
r4 2 32 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.0675 $X2=0.5005 $Y2=0.0675
r5 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0675 $X2=0.4860 $Y2=0.0675
r6 33 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4715 $Y2=0.0675
r7 3 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0675
+ $X2=0.5940 $Y2=0.0720
r8 2 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0675
+ $X2=0.4900 $Y2=0.0720
r9 28 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5805
+ $Y=0.0720 $X2=0.5940 $Y2=0.0720
r10 27 28 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0720 $X2=0.5805 $Y2=0.0720
r11 26 27 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.5420
+ $Y=0.0720 $X2=0.5670 $Y2=0.0720
r12 25 26 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5150
+ $Y=0.0720 $X2=0.5420 $Y2=0.0720
r13 24 25 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.4995
+ $Y=0.0720 $X2=0.5150 $Y2=0.0720
r14 23 24 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4900
+ $Y=0.0720 $X2=0.4995 $Y2=0.0720
r15 22 23 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4810
+ $Y=0.0720 $X2=0.4900 $Y2=0.0720
r16 21 22 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4620
+ $Y=0.0720 $X2=0.4810 $Y2=0.0720
r17 20 21 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4305
+ $Y=0.0720 $X2=0.4620 $Y2=0.0720
r18 19 20 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0720 $X2=0.4305 $Y2=0.0720
r19 18 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3915
+ $Y=0.0720 $X2=0.4050 $Y2=0.0720
r20 17 18 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0720 $X2=0.3915 $Y2=0.0720
r21 13 17 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3665
+ $Y=0.0720 $X2=0.3780 $Y2=0.0720
r22 1 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.0540
+ $X2=0.3780 $Y2=0.0720
r23 15 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r24 10 14 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3800 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r25 1 10 1e-05
.ends

.subckt PM_AO31x2_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00700704f
.ends

.subckt PM_AO31x2_ASAP7_75t_R%NET29 VSS 12 13 28 29 1 7 9 2 8
c1 1 VSS 0.00974681f
c2 2 VSS 0.00485877f
c3 7 VSS 0.00459825f
c4 8 VSS 0.00233864f
c5 9 VSS 0.0314344f
r1 29 27 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r2 2 27 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0675 $X2=0.4320 $Y2=0.0675
r4 28 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4175 $Y2=0.0675
r5 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4320 $Y2=0.0360
r6 23 24 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3935
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r7 22 23 13.6416 $w=1.3e-08 $l=5.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3350
+ $Y=0.0360 $X2=0.3935 $Y2=0.0360
r8 21 22 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.3350 $Y2=0.0360
r9 20 21 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.2970 $Y2=0.0360
r10 19 20 10.2603 $w=1.3e-08 $l=4.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2260
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r11 18 19 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1720
+ $Y=0.0360 $X2=0.2260 $Y2=0.0360
r12 17 18 9.67737 $w=1.3e-08 $l=4.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1305
+ $Y=0.0360 $X2=0.1720 $Y2=0.0360
r13 16 17 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1120
+ $Y=0.0360 $X2=0.1305 $Y2=0.0360
r14 14 16 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1030
+ $Y=0.0360 $X2=0.1120 $Y2=0.0360
r15 9 14 1.39914 $w=1.3e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.0970
+ $Y=0.0360 $X2=0.1030 $Y2=0.0360
r16 1 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1120 $Y2=0.0360
r17 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r18 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r19 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r20 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.0935 $Y2=0.0675
.ends

.subckt PM_AO31x2_ASAP7_75t_R%A3 VSS 21 3 4 7 1 10
c1 1 VSS 0.00880922f
c2 3 VSS 0.080456f
c3 4 VSS 0.0803375f
c4 5 VSS 0.0113851f
c5 6 VSS 0.00538462f
c6 7 VSS 0.00323729f
c7 8 VSS 0.00994999f
c8 9 VSS 0.00279821f
c9 10 VSS 0.00498239f
r1 8 27 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0360 $X2=0.0270 $Y2=0.0540
r2 6 9 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1665 $X2=0.0270 $Y2=0.1350
r3 6 10 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1665 $X2=0.0270 $Y2=0.1980
r4 26 27 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0720 $X2=0.0270 $Y2=0.0540
r5 5 9 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1035 $X2=0.0270 $Y2=0.1350
r6 5 26 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1035 $X2=0.0270 $Y2=0.0720
r7 9 23 3.60008 $w=1.51951e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1350 $X2=0.0475 $Y2=0.1350
r8 4 19 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r9 21 7 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0655 $Y2=0.1350
r10 7 23 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0655
+ $Y=0.1350 $X2=0.0475 $Y2=0.1350
r11 17 19 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1350 $X2=0.1350 $Y2=0.1350
r12 16 17 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1350 $X2=0.1225 $Y2=0.1350
r13 15 16 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1350 $X2=0.1080 $Y2=0.1350
r14 13 15 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0905 $Y=0.1350 $X2=0.0935 $Y2=0.1350
r15 12 13 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0905 $Y2=0.1350
r16 21 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
r17 1 12 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r18 1 14 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1350 $X2=0.0705 $Y2=0.1350
r19 3 12 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0810 $Y2=0.1350
r20 3 14 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.0810 $Y=0.1350 $X2=0.0705 $Y2=0.1350
r21 3 15 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1350
.ends

.subckt PM_AO31x2_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.004084f
.ends

.subckt PM_AO31x2_ASAP7_75t_R%NET23 VSS 23 26 43 45 48 49 52 53 1 16 2 17 21 3
+ 18 4 19 5 20
c1 1 VSS 0.00808224f
c2 2 VSS 0.0070848f
c3 3 VSS 0.00544565f
c4 4 VSS 0.00971263f
c5 5 VSS 0.00955762f
c6 16 VSS 0.00368874f
c7 17 VSS 0.00334971f
c8 18 VSS 0.00229114f
c9 19 VSS 0.00456086f
c10 20 VSS 0.0044963f
c11 21 VSS 0.0446677f
r1 53 51 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r2 5 51 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5400 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r3 20 5 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.2025 $X2=0.5400 $Y2=0.2025
r4 52 20 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.2025 $X2=0.5255 $Y2=0.2025
r5 49 47 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r6 4 47 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r7 19 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r8 48 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r9 18 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2680 $Y2=0.2025
r10 45 18 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r11 43 42 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r12 16 42 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r13 5 40 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.2025
+ $X2=0.5400 $Y2=0.2340
r14 4 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.2340
r15 3 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.2340
r16 1 31 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0520 $Y2=0.2340
r17 39 40 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.2340 $X2=0.5400 $Y2=0.2340
r18 38 39 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4860 $Y2=0.2340
r19 37 38 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.2340 $X2=0.4320 $Y2=0.2340
r20 36 37 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.3510 $Y2=0.2340
r21 35 36 9.32759 $w=1.3e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2300
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r22 34 35 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1850
+ $Y=0.2340 $X2=0.2300 $Y2=0.2340
r23 33 34 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1850 $Y2=0.2340
r24 32 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r25 28 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0610
+ $Y=0.2340 $X2=0.0790 $Y2=0.2340
r26 28 31 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0610
+ $Y=0.2340 $X2=0.0520 $Y2=0.2340
r27 27 29 5.13018 $w=1.3e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1010
+ $Y=0.2340 $X2=0.0790 $Y2=0.2340
r28 21 27 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1255
+ $Y=0.2340 $X2=0.1010 $Y2=0.2340
r29 21 32 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.1255
+ $Y=0.2340 $X2=0.1485 $Y2=0.2340
r30 2 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r31 26 25 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r32 24 25 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1720 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r33 2 24 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1600 $Y=0.2025 $X2=0.1720 $Y2=0.2025
r34 17 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1600 $Y2=0.2025
r35 23 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r36 1 16 1e-05
.ends

.subckt PM_AO31x2_ASAP7_75t_R%NET18 VSS 13 14 65 66 90 93 95 26 5 27 4 15 18 17
+ 19 28 24 20 6 23 16 31 30 32 1 25
c1 1 VSS 0.00889053f
c2 4 VSS 0.00560946f
c3 5 VSS 0.00296339f
c4 6 VSS 0.00463474f
c5 13 VSS 0.0814247f
c6 14 VSS 0.0807269f
c7 15 VSS 0.00484967f
c8 16 VSS 0.00437403f
c9 17 VSS 0.0044079f
c10 18 VSS 0.00120882f
c11 19 VSS 0.0103146f
c12 20 VSS 0.0136433f
c13 21 VSS 0.000946878f
c14 22 VSS 0.00416918f
c15 23 VSS 0.00406858f
c16 24 VSS 0.00422736f
c17 25 VSS 0.00354248f
c18 26 VSS 0.000828615f
c19 27 VSS 0.00112005f
c20 28 VSS 0.00110063f
c21 29 VSS 0.003088f
c22 30 VSS 0.00327781f
c23 31 VSS 0.000461783f
c24 32 VSS 0.00389158f
r1 15 4 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0540 $X2=0.2140 $Y2=0.0540
r2 95 15 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0540 $X2=0.2015 $Y2=0.0540
r3 4 86 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0540
+ $X2=0.2160 $Y2=0.0720
r4 93 92 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r5 91 92 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2260 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r6 5 91 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2140 $Y=0.2025 $X2=0.2260 $Y2=0.2025
r7 17 5 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2140 $Y2=0.2025
r8 90 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r9 86 87 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0720 $X2=0.2295 $Y2=0.0720
r10 27 84 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0720 $X2=0.2430 $Y2=0.1035
r11 27 87 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0720 $X2=0.2295 $Y2=0.0720
r12 5 78 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.1980
r13 83 84 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1035
r14 82 83 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1485 $X2=0.2430 $Y2=0.1350
r15 81 82 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1620 $X2=0.2430 $Y2=0.1485
r16 18 26 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1800 $X2=0.2430 $Y2=0.1980
r17 18 81 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1800 $X2=0.2430 $Y2=0.1620
r18 78 79 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1980 $X2=0.2295 $Y2=0.1980
r19 26 76 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.1980 $X2=0.2700 $Y2=0.1980
r20 26 79 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.1980 $X2=0.2295 $Y2=0.1980
r21 75 76 8.51143 $w=1.3e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.3065
+ $Y=0.1980 $X2=0.2700 $Y2=0.1980
r22 74 75 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3605
+ $Y=0.1980 $X2=0.3065 $Y2=0.1980
r23 73 74 10.3769 $w=1.3e-08 $l=4.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1980 $X2=0.3605 $Y2=0.1980
r24 72 73 10.3769 $w=1.3e-08 $l=4.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.4495
+ $Y=0.1980 $X2=0.4050 $Y2=0.1980
r25 71 72 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.5035
+ $Y=0.1980 $X2=0.4495 $Y2=0.1980
r26 70 71 8.04505 $w=1.3e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.5380
+ $Y=0.1980 $X2=0.5035 $Y2=0.1980
r27 69 70 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5560
+ $Y=0.1980 $X2=0.5380 $Y2=0.1980
r28 68 69 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1980 $X2=0.5560 $Y2=0.1980
r29 67 68 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.5920
+ $Y=0.1980 $X2=0.5670 $Y2=0.1980
r30 19 28 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6100 $Y=0.1980 $X2=0.6210 $Y2=0.1980
r31 19 67 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6100
+ $Y=0.1980 $X2=0.5920 $Y2=0.1980
r32 21 29 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.2160 $X2=0.6210 $Y2=0.2340
r33 21 28 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.2160 $X2=0.6210 $Y2=0.1980
r34 66 64 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.0675 $X2=0.5545 $Y2=0.0675
r35 6 64 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5400 $Y=0.0675 $X2=0.5545 $Y2=0.0675
r36 16 6 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.0675 $X2=0.5400 $Y2=0.0675
r37 65 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.0675 $X2=0.5255 $Y2=0.0675
r38 6 61 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.0675
+ $X2=0.5400 $Y2=0.0360
r39 22 32 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6480 $Y=0.2340 $X2=0.6750 $Y2=0.2340
r40 22 29 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6480 $Y=0.2340 $X2=0.6210 $Y2=0.2340
r41 61 62 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.0360 $X2=0.5785 $Y2=0.0360
r42 59 62 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.6190
+ $Y=0.0360 $X2=0.5785 $Y2=0.0360
r43 20 30 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6480 $Y=0.0360 $X2=0.6750 $Y2=0.0360
r44 20 59 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6480
+ $Y=0.0360 $X2=0.6190 $Y2=0.0360
r45 32 58 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6750 $Y=0.2340 $X2=0.6750 $Y2=0.2070
r46 30 54 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0360 $X2=0.6750 $Y2=0.0540
r47 57 58 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1800 $X2=0.6750 $Y2=0.2070
r48 56 57 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1620 $X2=0.6750 $Y2=0.1800
r49 55 56 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1510 $X2=0.6750 $Y2=0.1620
r50 24 31 1.50137 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6750 $Y=0.1465 $X2=0.6750 $Y2=0.1350
r51 24 55 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1465 $X2=0.6750 $Y2=0.1510
r52 53 54 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0720 $X2=0.6750 $Y2=0.0540
r53 52 53 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0900 $X2=0.6750 $Y2=0.0720
r54 23 31 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1125 $X2=0.6750 $Y2=0.1350
r55 23 52 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1125 $X2=0.6750 $Y2=0.0900
r56 14 42 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.7830 $Y=0.1350 $X2=0.7830 $Y2=0.1350
r57 48 49 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.7580
+ $Y=0.1350 $X2=0.7830 $Y2=0.1350
r58 47 48 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.7415
+ $Y=0.1350 $X2=0.7580 $Y2=0.1350
r59 46 47 0.46638 $w=1.3e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.7395
+ $Y=0.1350 $X2=0.7415 $Y2=0.1350
r60 45 46 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1350 $X2=0.7395 $Y2=0.1350
r61 25 45 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.1350 $X2=0.7290 $Y2=0.1350
r62 25 31 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7020 $Y=0.1350 $X2=0.6750 $Y2=0.1350
r63 42 49 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7830 $Y=0.1350
+ $X2=0.7830 $Y2=0.1350
r64 41 42 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.7735
+ $Y=0.1350 $X2=0.7830 $Y2=0.1350
r65 39 41 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.7705 $Y=0.1350 $X2=0.7735 $Y2=0.1350
r66 38 39 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7560 $Y=0.1350 $X2=0.7705 $Y2=0.1350
r67 37 38 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7415 $Y=0.1350 $X2=0.7560 $Y2=0.1350
r68 35 37 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.7385 $Y=0.1350 $X2=0.7415 $Y2=0.1350
r69 34 35 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.7290
+ $Y=0.1350 $X2=0.7385 $Y2=0.1350
r70 34 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7290 $Y=0.1350
+ $X2=0.7290 $Y2=0.1350
r71 1 34 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.7195
+ $Y=0.1350 $X2=0.7290 $Y2=0.1350
r72 1 36 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.7195
+ $Y=0.1350 $X2=0.7185 $Y2=0.1350
r73 13 34 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.7290 $Y=0.1350 $X2=0.7290 $Y2=0.1350
r74 13 36 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.7290 $Y=0.1350 $X2=0.7185 $Y2=0.1350
r75 13 37 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.7290 $Y=0.1350 $X2=0.7415 $Y2=0.1350
.ends

.subckt PM_AO31x2_ASAP7_75t_R%B VSS 21 3 4 8 5 6 10 7 1 9
c1 1 VSS 0.00760653f
c2 3 VSS 0.0445046f
c3 4 VSS 0.00785578f
c4 5 VSS 0.00298137f
c5 6 VSS 0.00281393f
c6 7 VSS 0.00281673f
c7 8 VSS 0.00319244f
c8 9 VSS 0.00334737f
c9 10 VSS 0.00217709f
r1 6 10 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1665 $X2=0.1350 $Y2=0.1350
r2 6 9 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1665 $X2=0.1350 $Y2=0.1980
r3 5 10 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1035 $X2=0.1350 $Y2=0.1350
r4 5 8 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1035 $X2=0.1350 $Y2=0.0720
r5 4 19 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r6 21 7 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1620 $Y2=0.1350
r7 7 10 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1620 $Y=0.1350 $X2=0.1350 $Y2=0.1350
r8 17 19 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2305 $Y=0.1350 $X2=0.2430 $Y2=0.1350
r9 16 17 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2160 $Y=0.1350 $X2=0.2305 $Y2=0.1350
r10 15 16 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2015 $Y=0.1350 $X2=0.2160 $Y2=0.1350
r11 13 15 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1985 $Y=0.1350 $X2=0.2015 $Y2=0.1350
r12 12 13 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1985 $Y2=0.1350
r13 21 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
r14 1 12 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1795
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r15 1 14 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.1795
+ $Y=0.1350 $X2=0.1785 $Y2=0.1350
r16 3 12 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1890 $Y2=0.1350
r17 3 14 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.1890 $Y=0.1350 $X2=0.1785 $Y2=0.1350
r18 3 15 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1890 $Y=0.1350 $X2=0.2015 $Y2=0.1350
.ends


*
.SUBCKT AO31x2_ASAP7_75t_R VSS VDD A3 B A2 A1 Y
*
* VSS VSS
* VDD VDD
* A3 A3
* B B
* A2 A2
* A1 A1
* Y Y
*
*

MM4 N_MM4_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@2 N_MM4@2_d N_MM10@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM9_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM7_g N_MM3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3@2 N_MM3@2_d N_MM7@2_g N_MM3@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM6_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2@2 N_MM2@2_d N_MM6@2_g N_MM2@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM1_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@2 N_MM0@2_d N_MM1@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10@2 N_MM10@2_d N_MM10@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9@2 N_MM9@2_d N_MM9@2_g N_MM9@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7@2 N_MM7@2_d N_MM7@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM6_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6@2 N_MM6@2_d N_MM6@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1@2 N_MM1@2_d N_MM1@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AO31x2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AO31x2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AO31x2_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_AO31x2_ASAP7_75t_R%noxref_13
cc_1 N_noxref_13_1 N_MM4_g 0.00220221f
cc_2 N_noxref_13_1 N_NET23_16 0.0359811f
cc_3 N_noxref_13_1 N_noxref_12_1 0.00176823f
x_PM_AO31x2_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_AO31x2_ASAP7_75t_R%noxref_17
cc_4 N_noxref_17_1 N_MM7_g 0.00160168f
cc_5 N_noxref_17_1 N_NET23_19 0.000666455f
cc_6 N_noxref_17_1 N_noxref_14_1 0.000477972f
cc_7 N_noxref_17_1 N_noxref_15_1 0.00766649f
cc_8 N_noxref_17_1 N_noxref_16_1 0.00123366f
x_PM_AO31x2_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_AO31x2_ASAP7_75t_R%noxref_12
cc_9 N_noxref_12_1 N_MM4_g 0.00227979f
cc_10 N_noxref_12_1 N_NET23_16 0.000476466f
x_PM_AO31x2_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_AO31x2_ASAP7_75t_R%noxref_19
cc_11 N_noxref_19_1 N_MM6@2_g 0.00141215f
cc_12 N_noxref_19_1 N_noxref_18_1 0.00123633f
x_PM_AO31x2_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_AO31x2_ASAP7_75t_R%noxref_21
cc_13 N_noxref_21_1 N_MM1_g 0.00178196f
cc_14 N_noxref_21_1 N_noxref_19_1 0.00766591f
cc_15 N_noxref_21_1 N_noxref_20_1 0.00123835f
x_PM_AO31x2_ASAP7_75t_R%Y VSS Y N_MM0_d N_MM0@2_d N_MM1_d N_MM1@2_d N_Y_7
+ N_Y_10 N_Y_8 N_Y_1 N_Y_11 N_Y_2 PM_AO31x2_ASAP7_75t_R%Y
cc_16 N_Y_7 N_NET18_30 0.000133584f
cc_17 N_Y_7 N_NET18_32 0.000170992f
cc_18 N_Y_7 N_NET18_24 0.000434808f
cc_19 N_Y_7 N_NET18_23 0.000451669f
cc_20 N_Y_7 N_NET18_1 0.000511993f
cc_21 N_Y_7 N_NET18_25 0.000743135f
cc_22 N_Y_10 N_NET18_25 0.000763846f
cc_23 N_Y_8 N_MM1@2_g 0.0307926f
cc_24 N_Y_1 N_NET18_1 0.000900397f
cc_25 N_Y_11 N_NET18_25 0.00191357f
cc_26 N_Y_1 N_MM1@2_g 0.00225164f
cc_27 N_Y_2 N_MM1@2_g 0.00227011f
cc_28 N_Y_1 N_NET18_25 0.00255298f
cc_29 N_Y_8 N_NET18_1 0.00418521f
cc_30 N_Y_7 N_MM1_g 0.0371983f
cc_31 N_Y_7 N_MM1@2_g 0.0685203f
x_PM_AO31x2_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_AO31x2_ASAP7_75t_R%noxref_23
cc_32 N_noxref_23_1 N_MM1@2_g 0.00150179f
cc_33 N_noxref_23_1 N_Y_8 0.00083234f
cc_34 N_noxref_23_1 N_noxref_22_1 0.0017734f
x_PM_AO31x2_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_AO31x2_ASAP7_75t_R%noxref_22
cc_35 N_noxref_22_1 N_MM1@2_g 0.00150086f
cc_36 N_noxref_22_1 N_Y_7 0.000827813f
x_PM_AO31x2_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_AO31x2_ASAP7_75t_R%noxref_16
cc_37 N_noxref_16_1 N_MM7_g 0.00171416f
cc_38 N_noxref_16_1 N_NET30_10 0.0356159f
cc_39 N_noxref_16_1 N_noxref_14_1 0.00784257f
x_PM_AO31x2_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_AO31x2_ASAP7_75t_R%noxref_18
cc_40 N_noxref_18_1 N_MM6@2_g 0.00142821f
cc_41 N_noxref_18_1 N_NET30_12 0.0354616f
x_PM_AO31x2_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_AO31x2_ASAP7_75t_R%noxref_20
cc_42 N_noxref_20_1 N_MM1_g 0.00174813f
cc_43 N_noxref_20_1 N_NET30_12 0.000566972f
cc_44 N_noxref_20_1 N_noxref_18_1 0.00766611f
x_PM_AO31x2_ASAP7_75t_R%A1 VSS A1 N_MM6_g N_MM6@2_g N_A1_9 N_A1_1 N_A1_7 N_A1_6
+ N_A1_8 PM_AO31x2_ASAP7_75t_R%A1
cc_45 N_MM6_g N_MM7@2_g 0.0055176f
x_PM_AO31x2_ASAP7_75t_R%A2 VSS A2 N_MM7_g N_MM7@2_g N_A2_9 N_A2_7 N_A2_5 N_A2_8
+ N_A2_1 N_A2_6 PM_AO31x2_ASAP7_75t_R%A2
x_PM_AO31x2_ASAP7_75t_R%NET30 VSS N_MM3_d N_MM3@2_d N_MM2_s N_MM2@2_s N_NET30_2
+ N_NET30_1 N_NET30_13 N_NET30_11 N_NET30_10 N_NET30_3 N_NET30_12
+ PM_AO31x2_ASAP7_75t_R%NET30
cc_46 N_NET30_2 N_MM7@2_g 0.000731282f
cc_47 N_NET30_1 N_MM7_g 0.00149849f
cc_48 N_NET30_13 N_A2_9 0.00156224f
cc_49 N_NET30_11 N_A2_1 0.00181007f
cc_50 N_NET30_13 N_A2_6 0.00218968f
cc_51 N_NET30_13 N_A2_1 0.00275287f
cc_52 N_NET30_11 N_MM7@2_g 0.0328291f
cc_53 N_NET30_10 N_MM7_g 0.035291f
cc_54 N_NET30_11 N_MM6@2_g 0.000435794f
cc_55 N_NET30_2 N_MM6_g 0.000952239f
cc_56 N_NET30_3 N_MM6@2_g 0.00106702f
cc_57 N_NET30_13 N_A1_6 0.00123115f
cc_58 N_NET30_13 N_A1_9 0.00135811f
cc_59 N_NET30_12 N_A1_1 0.00173939f
cc_60 N_NET30_13 N_A1_8 0.00487238f
cc_61 N_NET30_11 N_MM6_g 0.0329333f
cc_62 N_NET30_12 N_MM6@2_g 0.0348053f
cc_63 N_NET30_13 N_NET18_16 9.62401e-20
cc_64 N_NET30_13 N_NET18_24 0.000116348f
cc_65 N_NET30_13 N_NET18_31 0.000126716f
cc_66 N_NET30_13 N_NET18_6 0.00114792f
cc_67 N_NET30_13 N_NET18_19 0.000295888f
cc_68 N_NET30_13 N_NET18_23 0.000525299f
cc_69 N_NET30_11 N_NET18_16 0.000556225f
cc_70 N_NET30_3 N_NET18_20 0.000592472f
cc_71 N_NET30_12 N_NET18_16 0.00175846f
cc_72 N_NET30_2 N_NET18_6 0.00124509f
cc_73 N_NET30_3 N_NET18_6 0.00497004f
cc_74 N_NET30_13 N_NET18_20 0.00936799f
cc_75 N_NET30_10 N_NET29_8 0.000596655f
cc_76 N_NET30_13 N_NET29_2 0.000865916f
cc_77 N_NET30_11 N_NET29_8 0.00111854f
cc_78 N_NET30_1 N_NET29_2 0.00173545f
cc_79 N_NET30_2 N_NET29_2 0.00430519f
cc_80 N_NET30_13 N_NET29_9 0.0101749f
x_PM_AO31x2_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_AO31x2_ASAP7_75t_R%noxref_15
cc_81 N_noxref_15_1 N_MM9@2_g 0.00152878f
cc_82 N_noxref_15_1 N_NET23_18 0.0358316f
cc_83 N_noxref_15_1 N_noxref_14_1 0.00137221f
x_PM_AO31x2_ASAP7_75t_R%NET29 VSS N_MM4_d N_MM4@2_d N_MM3_s N_MM3@2_s N_NET29_1
+ N_NET29_7 N_NET29_9 N_NET29_2 N_NET29_8 PM_AO31x2_ASAP7_75t_R%NET29
cc_84 N_NET29_1 N_MM10@2_g 0.00198486f
cc_85 N_NET29_7 N_A3_1 0.00205218f
cc_86 N_NET29_7 N_MM4_g 0.0183374f
cc_87 N_NET29_7 N_MM10@2_g 0.0506657f
cc_88 N_NET29_9 N_B_8 0.00230193f
cc_89 N_NET29_9 N_MM9@2_g 0.00432803f
cc_90 N_NET29_2 N_MM7@2_g 0.00194522f
cc_91 N_NET29_8 N_A2_1 0.00222791f
cc_92 N_NET29_9 N_A2_7 0.00296852f
cc_93 N_NET29_8 N_MM7_g 0.0183444f
cc_94 N_NET29_8 N_MM7@2_g 0.0500456f
cc_95 N_NET29_9 N_NET18_18 0.000265635f
cc_96 N_NET29_9 N_NET18_4 0.000906422f
cc_97 N_NET29_9 N_NET18_27 0.00668737f
x_PM_AO31x2_ASAP7_75t_R%A3 VSS A3 N_MM4_g N_MM10@2_g N_A3_7 N_A3_1 N_A3_10
+ PM_AO31x2_ASAP7_75t_R%A3
x_PM_AO31x2_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_AO31x2_ASAP7_75t_R%noxref_14
cc_98 N_noxref_14_1 N_MM9@2_g 0.00888825f
cc_99 N_noxref_14_1 N_MM7_g 0.000738075f
cc_100 N_noxref_14_1 N_NET18_15 0.000751253f
cc_101 N_noxref_14_1 N_NET23_18 0.000504726f
cc_102 N_noxref_14_1 N_NET29_9 0.000307007f
cc_103 N_noxref_14_1 N_NET30_10 0.000625067f
x_PM_AO31x2_ASAP7_75t_R%NET23 VSS N_MM10@2_d N_MM9_s N_MM10_d N_MM9@2_s N_MM7_d
+ N_MM7@2_d N_MM6_d N_MM6@2_d N_NET23_1 N_NET23_16 N_NET23_2 N_NET23_17
+ N_NET23_21 N_NET23_3 N_NET23_18 N_NET23_4 N_NET23_19 N_NET23_5 N_NET23_20
+ PM_AO31x2_ASAP7_75t_R%NET23
cc_104 N_NET23_1 N_MM10@2_g 0.00130528f
cc_105 N_NET23_16 N_MM10@2_g 0.00048996f
cc_106 N_NET23_2 N_MM10@2_g 0.000704854f
cc_107 N_NET23_17 N_A3_1 0.00155516f
cc_108 N_NET23_21 N_MM10@2_g 0.00160243f
cc_109 N_NET23_21 N_A3_10 0.00195284f
cc_110 N_NET23_1 N_MM4_g 0.00202943f
cc_111 N_NET23_16 N_MM4_g 0.0333018f
cc_112 N_NET23_17 N_MM10@2_g 0.0341626f
cc_113 N_NET23_2 N_MM9@2_g 0.000817876f
cc_114 N_NET23_17 N_MM9@2_g 0.000394238f
cc_115 N_NET23_3 N_MM9@2_g 0.000821723f
cc_116 N_NET23_2 N_MM9_g 0.00147295f
cc_117 N_NET23_18 N_B_1 0.00171848f
cc_118 N_NET23_21 N_B_9 0.00227347f
cc_119 N_NET23_21 N_MM9@2_g 0.0023832f
cc_120 N_NET23_17 N_MM9_g 0.0330782f
cc_121 N_NET23_18 N_MM9@2_g 0.0347306f
cc_122 N_NET23_4 N_MM7@2_g 0.00210796f
cc_123 N_NET23_21 N_MM7@2_g 0.000302445f
cc_124 N_NET23_3 N_MM7@2_g 0.000774008f
cc_125 N_NET23_19 N_A2_1 0.0020607f
cc_126 N_NET23_19 N_MM7_g 0.0183278f
cc_127 N_NET23_19 N_MM7@2_g 0.0495957f
cc_128 N_NET23_5 N_MM6@2_g 0.00229458f
cc_129 N_NET23_20 N_A1_1 0.00201963f
cc_130 N_NET23_20 N_MM6_g 0.0183384f
cc_131 N_NET23_20 N_MM6@2_g 0.0496337f
cc_132 N_NET23_21 N_NET18_17 9.8447e-20
cc_133 N_NET23_21 N_NET18_5 0.000939909f
cc_134 N_NET23_4 N_NET18_19 0.00119429f
cc_135 N_NET23_3 N_NET18_18 0.000485623f
cc_136 N_NET23_5 N_NET18_19 0.00124274f
cc_137 N_NET23_17 N_NET18_17 0.000560377f
cc_138 N_NET23_3 N_NET18_19 0.000610518f
cc_139 N_NET23_18 N_NET18_17 0.00174244f
cc_140 N_NET23_2 N_NET18_5 0.00138013f
cc_141 N_NET23_21 N_NET18_26 0.00245379f
cc_142 N_NET23_3 N_NET18_5 0.00504124f
cc_143 N_NET23_21 N_NET18_19 0.0271202f
x_PM_AO31x2_ASAP7_75t_R%NET18 VSS N_MM1_g N_MM1@2_g N_MM2_d N_MM2@2_d N_MM9_d
+ N_MM9@2_d N_MM5_d N_NET18_26 N_NET18_5 N_NET18_27 N_NET18_4 N_NET18_15
+ N_NET18_18 N_NET18_17 N_NET18_19 N_NET18_28 N_NET18_24 N_NET18_20 N_NET18_6
+ N_NET18_23 N_NET18_16 N_NET18_31 N_NET18_30 N_NET18_32 N_NET18_1 N_NET18_25
+ PM_AO31x2_ASAP7_75t_R%NET18
cc_144 N_NET18_26 N_MM9@2_g 0.000428015f
cc_145 N_NET18_5 N_MM9@2_g 0.00275487f
cc_146 N_NET18_27 N_MM9@2_g 0.000205017f
cc_147 N_NET18_4 N_MM9@2_g 0.00143131f
cc_148 N_NET18_27 N_B_7 0.000698019f
cc_149 N_NET18_15 N_MM9_g 0.00892878f
cc_150 N_NET18_18 N_B_7 0.002018f
cc_151 N_NET18_26 N_B_7 0.00219693f
cc_152 N_NET18_17 N_B_1 0.00398608f
cc_153 N_NET18_15 N_MM9@2_g 0.0150504f
cc_154 N_NET18_17 N_MM9_g 0.0325947f
cc_155 N_NET18_17 N_MM9@2_g 0.0649808f
cc_156 N_NET18_27 N_A2_9 0.000374127f
cc_157 N_NET18_18 N_A2_7 0.00136177f
cc_158 N_NET18_18 N_A2_5 0.002778f
cc_159 N_NET18_19 N_A2_8 0.00283333f
cc_160 N_NET18_19 N_A2_9 0.00600333f
cc_161 N_NET18_28 N_MM6@2_g 0.000152975f
cc_162 N_NET18_24 N_MM6@2_g 0.000154056f
cc_163 N_NET18_20 N_MM6@2_g 0.000170572f
cc_164 N_NET18_6 N_MM6@2_g 0.00349186f
cc_165 N_NET18_23 N_MM6@2_g 0.000204972f
cc_166 N_NET18_19 N_MM6@2_g 0.000376825f
cc_167 N_NET18_19 N_A1_9 0.0010433f
cc_168 N_NET18_16 N_A1_1 0.00238925f
cc_169 N_NET18_19 N_A1_7 0.00561774f
cc_170 N_NET18_16 N_MM6_g 0.0189539f
cc_171 N_NET18_16 N_MM6@2_g 0.0509334f
x_PM_AO31x2_ASAP7_75t_R%B VSS B N_MM9_g N_MM9@2_g N_B_8 N_B_5 N_B_6 N_B_10
+ N_B_7 N_B_1 N_B_9 PM_AO31x2_ASAP7_75t_R%B
cc_172 N_B_8 N_MM10@2_g 0.000559567f
cc_173 N_B_5 N_A3_7 0.000692152f
cc_174 N_B_6 N_A3_7 0.000720854f
cc_175 N_B_10 N_A3_1 0.00127367f
cc_176 N_B_10 N_A3_7 0.00186843f
cc_177 N_MM9_g N_MM10@2_g 0.00590746f
*END of AO31x2_ASAP7_75t_R.pxi
.ENDS
** Design:	AO322x2_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AO322x2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AO322x2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AO322x2_ASAP7_75t_R%NET50 VSS 2 3 1
c1 1 VSS 0.000851044f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0540 $X2=0.4860 $Y2=0.0540
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0540 $X2=0.4860 $Y2=0.0540
.ends

.subckt PM_AO322x2_ASAP7_75t_R%NET52 VSS 2 3 1
c1 1 VSS 0.000960467f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_AO322x2_ASAP7_75t_R%NET49 VSS 2 3 1
c1 1 VSS 0.000961232f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_AO322x2_ASAP7_75t_R%NET51 VSS 2 3 1
c1 1 VSS 0.000884641f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0540 $X2=0.2700 $Y2=0.0540
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0540 $X2=0.2700 $Y2=0.0540
.ends

.subckt PM_AO322x2_ASAP7_75t_R%NET27 VSS 20 21 37 40 42 10 13 1 16 11 2 15 12 3
c1 1 VSS 0.00953298f
c2 2 VSS 0.0057054f
c3 3 VSS 0.00433309f
c4 10 VSS 0.00453792f
c5 11 VSS 0.00330406f
c6 12 VSS 0.00271266f
c7 13 VSS 0.00850305f
c8 14 VSS 0.000585153f
c9 15 VSS 0.00211261f
c10 16 VSS 0.000587655f
c11 17 VSS 0.00309278f
r1 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3220 $Y2=0.2025
r2 42 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r3 40 39 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r4 38 39 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2260 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r5 2 38 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2140 $Y=0.2025 $X2=0.2260 $Y2=0.2025
r6 11 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2140 $Y2=0.2025
r7 37 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r8 3 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3200 $Y2=0.1980
r9 2 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.1980
r10 32 33 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3015
+ $Y=0.1980 $X2=0.3200 $Y2=0.1980
r11 31 32 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2720
+ $Y=0.1980 $X2=0.3015 $Y2=0.1980
r12 30 31 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2540
+ $Y=0.1980 $X2=0.2720 $Y2=0.1980
r13 29 30 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1980 $X2=0.2540 $Y2=0.1980
r14 28 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.1980 $X2=0.2430 $Y2=0.1980
r15 27 28 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1980 $X2=0.2295 $Y2=0.1980
r16 15 27 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2025
+ $Y=0.1980 $X2=0.2160 $Y2=0.1980
r17 15 16 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2025 $Y=0.1980 $X2=0.1890 $Y2=0.1980
r18 14 17 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2160 $X2=0.1890 $Y2=0.2340
r19 14 16 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2160 $X2=0.1890 $Y2=0.1980
r20 17 26 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2340 $X2=0.1620 $Y2=0.2340
r21 25 26 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1305
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r22 24 25 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1120
+ $Y=0.2340 $X2=0.1305 $Y2=0.2340
r23 22 24 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1030
+ $Y=0.2340 $X2=0.1120 $Y2=0.2340
r24 13 22 1.39914 $w=1.3e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.0970
+ $Y=0.2340 $X2=0.1030 $Y2=0.2340
r25 1 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1120 $Y2=0.2340
r26 20 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r27 1 19 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r28 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r29 21 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
.ends

.subckt PM_AO322x2_ASAP7_75t_R%A3 VSS 6 3 1 4
c1 1 VSS 0.00742725f
c2 3 VSS 0.083401f
c3 4 VSS 0.0040853f
r1 7 8 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1085 $X2=0.1890 $Y2=0.1350
r2 6 7 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0905 $X2=0.1890 $Y2=0.1085
r3 6 4 1.16595 $w=1.3e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0905 $X2=0.1890 $Y2=0.0855
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AO322x2_ASAP7_75t_R%B2 VSS 8 3 1 4
c1 1 VSS 0.00749328f
c2 3 VSS 0.0466616f
c3 4 VSS 0.00487207f
r1 8 7 0.816164 $w=1.3e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1505 $X2=0.2430 $Y2=0.1470
r2 6 7 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1470
r3 4 6 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1035 $X2=0.2430 $Y2=0.1350
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r5 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AO322x2_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.00523085f
.ends

.subckt PM_AO322x2_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.0419678f
.ends

.subckt PM_AO322x2_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.00404866f
.ends

.subckt PM_AO322x2_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.00421494f
.ends

.subckt PM_AO322x2_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.00439679f
.ends

.subckt PM_AO322x2_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.0310996f
.ends

.subckt PM_AO322x2_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.00590787f
.ends

.subckt PM_AO322x2_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.00473718f
.ends

.subckt PM_AO322x2_ASAP7_75t_R%C1 VSS 6 3 1 4
c1 1 VSS 0.00639913f
c2 3 VSS 0.00877098f
c3 4 VSS 0.00463283f
r1 7 8 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1045 $X2=0.4590 $Y2=0.1350
r2 6 7 5.13018 $w=1.3e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0825 $X2=0.4590 $Y2=0.1045
r3 6 4 0.23319 $w=1.3e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0825 $X2=0.4590 $Y2=0.0815
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1350
+ $X2=0.4590 $Y2=0.1350
.ends

.subckt PM_AO322x2_ASAP7_75t_R%noxref_26 VSS 1
c1 1 VSS 0.00553129f
.ends

.subckt PM_AO322x2_ASAP7_75t_R%A2 VSS 13 3 6 5 1 4
c1 1 VSS 0.00505843f
c2 3 VSS 0.0458018f
c3 4 VSS 0.00324568f
c4 5 VSS 0.002276f
c5 6 VSS 0.00264415f
r1 13 6 0.510222 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1355
+ $Y=0.1980 $X2=0.1305 $Y2=0.1980
r2 5 8 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.0720 $X2=0.1350 $Y2=0.1035
r3 13 11 2.14973 $w=1.32632e-08 $l=1.80069e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1355 $Y=0.1980 $X2=0.1350 $Y2=0.1800
r4 10 11 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1675 $X2=0.1350 $Y2=0.1800
r5 9 10 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1540 $X2=0.1350 $Y2=0.1675
r6 4 8 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1035
r7 4 9 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1540
r8 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r9 1 4 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AO322x2_ASAP7_75t_R%C2 VSS 9 3 1 4 5
c1 1 VSS 0.00485283f
c2 3 VSS 0.0352783f
c3 4 VSS 0.00340993f
c4 5 VSS 0.00564301f
r1 9 8 0.932759 $w=1.3e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1515 $X2=0.5130 $Y2=0.1475
r2 7 8 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1475
r3 4 7 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1035 $X2=0.5130 $Y2=0.1350
r4 4 5 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1035 $X2=0.5130 $Y2=0.0720
r5 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r6 1 7 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.1350
+ $X2=0.5130 $Y2=0.1350
.ends

.subckt PM_AO322x2_ASAP7_75t_R%A1 VSS 14 3 6 1 4 7 9
c1 1 VSS 0.00246939f
c2 3 VSS 0.04324f
c3 4 VSS 0.00387183f
c4 5 VSS 0.00856242f
c5 6 VSS 0.00241454f
c6 7 VSS 0.00309219f
c7 8 VSS 0.00197799f
c8 9 VSS 0.00856174f
r1 9 18 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.2340 $X2=0.0270 $Y2=0.2160
r2 17 18 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1980 $X2=0.0270 $Y2=0.2160
r3 5 8 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1665 $X2=0.0270 $Y2=0.1350
r4 5 17 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1665 $X2=0.0270 $Y2=0.1980
r5 4 8 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1035 $X2=0.0270 $Y2=0.1350
r6 4 7 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1035 $X2=0.0270 $Y2=0.0720
r7 8 13 2.55073 $w=1.58125e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1350 $X2=0.0430 $Y2=0.1350
r8 14 15 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0505
+ $Y=0.1350 $X2=0.0530 $Y2=0.1350
r9 14 13 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0505
+ $Y=0.1350 $X2=0.0430 $Y2=0.1350
r10 6 11 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.0635
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r11 6 15 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0635
+ $Y=0.1350 $X2=0.0530 $Y2=0.1350
r12 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r13 1 11 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AO322x2_ASAP7_75t_R%noxref_27 VSS 1
c1 1 VSS 0.00454876f
.ends

.subckt PM_AO322x2_ASAP7_75t_R%noxref_29 VSS 1
c1 1 VSS 0.00518025f
.ends

.subckt PM_AO322x2_ASAP7_75t_R%B1 VSS 8 3 1 4 5 6
c1 1 VSS 0.00524318f
c2 3 VSS 0.00819523f
c3 4 VSS 0.00324629f
c4 5 VSS 0.00318719f
c5 6 VSS 0.00286065f
r1 6 11 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1620 $X2=0.2970 $Y2=0.1485
r2 10 11 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1485
r3 9 10 6.64591 $w=1.3e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1065 $X2=0.2970 $Y2=0.1350
r4 8 9 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0865 $X2=0.2970 $Y2=0.1065
r5 8 4 0.699569 $w=1.3e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0865 $X2=0.2970 $Y2=0.0835
r6 4 5 1.50137 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0835 $X2=0.2970 $Y2=0.0720
r7 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r8 1 10 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_AO322x2_ASAP7_75t_R%noxref_28 VSS 1
c1 1 VSS 0.00487665f
.ends

.subckt PM_AO322x2_ASAP7_75t_R%NET53 VSS 12 13 22 23 7 1 8 2 9
c1 1 VSS 0.0045545f
c2 2 VSS 0.00435935f
c3 7 VSS 0.00220815f
c4 8 VSS 0.00219336f
c5 9 VSS 0.0229228f
r1 23 21 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r2 2 21 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4860 $Y2=0.2025
r4 22 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r5 2 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2025
+ $X2=0.4860 $Y2=0.2340
r6 17 18 11.5429 $w=1.3e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4365
+ $Y=0.2340 $X2=0.4860 $Y2=0.2340
r7 16 17 16.2067 $w=1.3e-08 $l=6.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.3670
+ $Y=0.2340 $X2=0.4365 $Y2=0.2340
r8 15 16 13.6416 $w=1.3e-08 $l=5.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3085
+ $Y=0.2340 $X2=0.3670 $Y2=0.2340
r9 14 15 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.3085 $Y2=0.2340
r10 9 14 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2585
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r11 1 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.2340
r12 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r13 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r14 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r15 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
.ends

.subckt PM_AO322x2_ASAP7_75t_R%Y VSS 32 23 38 45 47 14 18 2 16 13 15 1 17 3 4 19
c1 1 VSS 0.00919811f
c2 2 VSS 0.00806027f
c3 3 VSS 0.00784251f
c4 4 VSS 0.00787568f
c5 13 VSS 0.00356745f
c6 14 VSS 0.00350409f
c7 15 VSS 0.00357196f
c8 16 VSS 0.00345596f
c9 17 VSS 0.0147747f
c10 18 VSS 0.0139694f
c11 19 VSS 0.00322547f
c12 20 VSS 0.00281433f
c13 21 VSS 0.00306474f
r1 47 46 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.2025 $X2=0.6625 $Y2=0.2025
r2 15 46 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6500 $Y=0.2025 $X2=0.6625 $Y2=0.2025
r3 16 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7415 $Y=0.2025 $X2=0.7540 $Y2=0.2025
r4 45 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.2025 $X2=0.7415 $Y2=0.2025
r5 2 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.2025
+ $X2=0.6480 $Y2=0.2340
r6 4 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7560 $Y=0.2025
+ $X2=0.7560 $Y2=0.2340
r7 42 43 12.1259 $w=1.3e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6480
+ $Y=0.2340 $X2=0.7000 $Y2=0.2340
r8 39 40 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.2340 $X2=0.7695 $Y2=0.2340
r9 18 39 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.7450
+ $Y=0.2340 $X2=0.7560 $Y2=0.2340
r10 18 43 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.7450
+ $Y=0.2340 $X2=0.7000 $Y2=0.2340
r11 21 36 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.2340 $X2=0.7830 $Y2=0.2160
r12 21 40 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7830 $Y=0.2340 $X2=0.7695 $Y2=0.2340
r13 14 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7415 $Y=0.0675 $X2=0.7540 $Y2=0.0675
r14 38 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.0675 $X2=0.7415 $Y2=0.0675
r15 35 36 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1755 $X2=0.7830 $Y2=0.2160
r16 34 35 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1350 $X2=0.7830 $Y2=0.1755
r17 33 34 3.38125 $w=1.3e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1205 $X2=0.7830 $Y2=0.1350
r18 32 33 1.39914 $w=1.3e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1145 $X2=0.7830 $Y2=0.1205
r19 32 31 3.96423 $w=1.3e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.1145 $X2=0.7830 $Y2=0.0975
r20 30 31 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.0720 $X2=0.7830 $Y2=0.0975
r21 19 20 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.0540 $X2=0.7830 $Y2=0.0360
r22 19 30 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7830
+ $Y=0.0540 $X2=0.7830 $Y2=0.0720
r23 3 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7560 $Y=0.0675
+ $X2=0.7560 $Y2=0.0360
r24 20 29 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7830 $Y=0.0360 $X2=0.7695 $Y2=0.0360
r25 28 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.0360 $X2=0.7695 $Y2=0.0360
r26 27 28 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.7450
+ $Y=0.0360 $X2=0.7560 $Y2=0.0360
r27 26 27 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.7000
+ $Y=0.0360 $X2=0.7450 $Y2=0.0360
r28 25 26 12.1259 $w=1.3e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6480
+ $Y=0.0360 $X2=0.7000 $Y2=0.0360
r29 17 25 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6365
+ $Y=0.0360 $X2=0.6480 $Y2=0.0360
r30 1 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.0540
+ $X2=0.6480 $Y2=0.0360
r31 23 22 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.0675 $X2=0.6625 $Y2=0.0675
r32 13 22 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6500 $Y=0.0675 $X2=0.6625 $Y2=0.0675
r33 2 15 1e-05
r34 1 13 1e-05
.ends

.subckt PM_AO322x2_ASAP7_75t_R%NET25 VSS 19 20 66 74 94 96 98 4 21 26 5 22 32
+ 27 7 6 23 31 28 24 8 30 33 29 25 34 1
c1 1 VSS 0.00982309f
c2 4 VSS 0.00660911f
c3 5 VSS 0.00529295f
c4 6 VSS 0.00608657f
c5 7 VSS 0.00365322f
c6 8 VSS 0.00404862f
c7 19 VSS 0.080229f
c8 20 VSS 0.0799626f
c9 21 VSS 0.00434562f
c10 22 VSS 0.00356841f
c11 23 VSS 0.00360877f
c12 24 VSS 0.0037617f
c13 25 VSS 0.00358288f
c14 26 VSS 0.033976f
c15 27 VSS 0.00234001f
c16 28 VSS 0.0024149f
c17 29 VSS 0.000877341f
c18 30 VSS 0.00428267f
c19 31 VSS 0.00630082f
c20 32 VSS 0.00136694f
c21 33 VSS 0.000523689f
c22 34 VSS 0.00117161f
r1 98 97 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r2 21 97 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r3 22 5 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0540 $X2=0.3220 $Y2=0.0540
r4 96 22 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0540 $X2=0.3095 $Y2=0.0540
r5 94 93 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0540 $X2=0.4465 $Y2=0.0540
r6 23 93 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4340 $Y=0.0540 $X2=0.4465 $Y2=0.0540
r7 4 92 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0500 $Y2=0.0360
r8 5 81 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0540
+ $X2=0.3200 $Y2=0.0360
r9 6 76 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0540
+ $X2=0.4320 $Y2=0.0360
r10 89 90 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0590
+ $Y=0.0360 $X2=0.0790 $Y2=0.0360
r11 89 92 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0590
+ $Y=0.0360 $X2=0.0500 $Y2=0.0360
r12 88 90 5.13017 $w=1.3e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1010
+ $Y=0.0360 $X2=0.0790 $Y2=0.0360
r13 87 88 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1255
+ $Y=0.0360 $X2=0.1010 $Y2=0.0360
r14 86 87 8.51143 $w=1.3e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1255 $Y2=0.0360
r15 85 86 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r16 84 85 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r17 83 84 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r18 82 83 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r19 80 81 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3015
+ $Y=0.0360 $X2=0.3200 $Y2=0.0360
r20 80 82 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3015
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r21 78 79 1.51573 $w=1.3e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3290
+ $Y=0.0360 $X2=0.3355 $Y2=0.0360
r22 78 81 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3290
+ $Y=0.0360 $X2=0.3200 $Y2=0.0360
r23 26 31 7.6809 $w=1.41842e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3670 $Y=0.0360 $X2=0.4050 $Y2=0.0360
r24 26 79 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3670
+ $Y=0.0360 $X2=0.3355 $Y2=0.0360
r25 75 76 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4185
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r26 31 72 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0360 $X2=0.4050 $Y2=0.0540
r27 31 75 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.0360 $X2=0.4185 $Y2=0.0360
r28 74 73 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r29 24 73 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4340 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r30 71 72 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0665 $X2=0.4050 $Y2=0.0540
r31 70 71 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0755 $X2=0.4050 $Y2=0.0665
r32 69 70 9.67738 $w=1.3e-08 $l=4.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1170 $X2=0.4050 $Y2=0.0755
r33 68 69 9.67738 $w=1.3e-08 $l=4.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1585 $X2=0.4050 $Y2=0.1170
r34 67 68 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1675 $X2=0.4050 $Y2=0.1585
r35 27 32 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1800 $X2=0.4050 $Y2=0.1980
r36 27 67 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1800 $X2=0.4050 $Y2=0.1675
r37 25 8 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.2025 $X2=0.5380 $Y2=0.2025
r38 66 25 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.2025 $X2=0.5255 $Y2=0.2025
r39 7 63 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4330 $Y2=0.1980
r40 32 62 1.61554 $w=1.62143e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.1980 $X2=0.4190 $Y2=0.1980
r41 8 56 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.2025
+ $X2=0.5360 $Y2=0.1980
r42 63 64 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4330
+ $Y=0.1980 $X2=0.4440 $Y2=0.1980
r43 62 63 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.4190
+ $Y=0.1980 $X2=0.4330 $Y2=0.1980
r44 61 64 0.932759 $w=1.3e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.4480
+ $Y=0.1980 $X2=0.4440 $Y2=0.1980
r45 60 61 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1980 $X2=0.4480 $Y2=0.1980
r46 59 60 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4840
+ $Y=0.1980 $X2=0.4590 $Y2=0.1980
r47 58 59 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5020
+ $Y=0.1980 $X2=0.4840 $Y2=0.1980
r48 57 58 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1980 $X2=0.5020 $Y2=0.1980
r49 55 56 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.5265
+ $Y=0.1980 $X2=0.5360 $Y2=0.1980
r50 55 57 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5265
+ $Y=0.1980 $X2=0.5130 $Y2=0.1980
r51 28 54 1.98211 $w=1.3e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.5450
+ $Y=0.1980 $X2=0.5535 $Y2=0.1980
r52 28 56 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5450
+ $Y=0.1980 $X2=0.5360 $Y2=0.1980
r53 34 53 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.1980 $X2=0.5670 $Y2=0.1765
r54 34 54 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.1980 $X2=0.5535 $Y2=0.1980
r55 29 33 2.78149 $w=1.76421e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.1540 $X2=0.5670 $Y2=0.1350
r56 29 53 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1540 $X2=0.5670 $Y2=0.1765
r57 20 44 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.7290 $Y=0.1350 $X2=0.7290 $Y2=0.1350
r58 49 50 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.1350 $X2=0.7290 $Y2=0.1350
r59 48 49 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1350 $X2=0.7020 $Y2=0.1350
r60 47 48 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.6500
+ $Y=0.1350 $X2=0.6750 $Y2=0.1350
r61 30 47 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.6050
+ $Y=0.1350 $X2=0.6500 $Y2=0.1350
r62 30 33 7.2121 $w=1.41842e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6050 $Y=0.1350 $X2=0.5670 $Y2=0.1350
r63 44 50 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7290 $Y=0.1350
+ $X2=0.7290 $Y2=0.1350
r64 43 44 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.7195
+ $Y=0.1350 $X2=0.7290 $Y2=0.1350
r65 41 43 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.7165 $Y=0.1350 $X2=0.7195 $Y2=0.1350
r66 40 41 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7020 $Y=0.1350 $X2=0.7165 $Y2=0.1350
r67 39 40 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6875 $Y=0.1350 $X2=0.7020 $Y2=0.1350
r68 37 39 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.6845 $Y=0.1350 $X2=0.6875 $Y2=0.1350
r69 36 37 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.6750
+ $Y=0.1350 $X2=0.6845 $Y2=0.1350
r70 36 48 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6750 $Y=0.1350
+ $X2=0.6750 $Y2=0.1350
r71 1 36 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.6655
+ $Y=0.1350 $X2=0.6750 $Y2=0.1350
r72 1 38 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.6655
+ $Y=0.1350 $X2=0.6645 $Y2=0.1350
r73 19 36 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.6750 $Y=0.1350 $X2=0.6750 $Y2=0.1350
r74 19 38 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.6750 $Y=0.1350 $X2=0.6645 $Y2=0.1350
r75 19 39 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.6750 $Y=0.1350 $X2=0.6875 $Y2=0.1350
r76 4 21 1e-05
r77 6 23 1e-05
r78 7 24 1e-05
.ends


*
.SUBCKT AO322x2_ASAP7_75t_R VSS VDD A1 A2 A3 B2 B1 C1 C2 Y
*
* VSS VSS
* VDD VDD
* A1 A1
* A2 A2
* A3 A3
* B2 B2
* B1 B1
* C1 C1
* C2 C2
* Y Y
*
*

MM0 N_MM0_d N_MM0_g N_MM0_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM10_g N_MM1_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM13_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM8_g N_MM3_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM9_g N_MM5_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM6 N_MM6_d N_MM12_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM16 N_MM16_d N_MM17_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM16@2 N_MM16@2_d N_MM17@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM13 N_MM13_d N_MM13_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 N_MM11_d N_MM11_g N_MM11_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM8_g N_MM8_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM12 N_MM12_d N_MM12_g N_MM12_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM17 N_MM17_d N_MM17_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM17@2 N_MM17@2_d N_MM17@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AO322x2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AO322x2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AO322x2_ASAP7_75t_R%NET50 VSS N_MM5_s N_MM6_d N_NET50_1
+ PM_AO322x2_ASAP7_75t_R%NET50
cc_1 N_NET50_1 N_MM9_g 0.0125302f
cc_2 N_NET50_1 N_MM12_g 0.0125382f
x_PM_AO322x2_ASAP7_75t_R%NET52 VSS N_MM1_s N_MM2_d N_NET52_1
+ PM_AO322x2_ASAP7_75t_R%NET52
cc_3 N_NET52_1 N_MM10_g 0.0173363f
cc_4 N_NET52_1 N_MM13_g 0.0173632f
x_PM_AO322x2_ASAP7_75t_R%NET49 VSS N_MM0_s N_MM1_d N_NET49_1
+ PM_AO322x2_ASAP7_75t_R%NET49
cc_5 N_NET49_1 N_MM0_g 0.0173236f
cc_6 N_NET49_1 N_MM10_g 0.0174877f
x_PM_AO322x2_ASAP7_75t_R%NET51 VSS N_MM4_d N_MM3_s N_NET51_1
+ PM_AO322x2_ASAP7_75t_R%NET51
cc_7 N_NET51_1 N_MM11_g 0.0126522f
cc_8 N_NET51_1 N_MM8_g 0.0127322f
x_PM_AO322x2_ASAP7_75t_R%NET27 VSS N_MM10_d N_MM7_d N_MM13_d N_MM11_s N_MM8_s
+ N_NET27_10 N_NET27_13 N_NET27_1 N_NET27_16 N_NET27_11 N_NET27_2 N_NET27_15
+ N_NET27_12 N_NET27_3 PM_AO322x2_ASAP7_75t_R%NET27
cc_9 N_NET27_10 N_A1_1 0.00077733f
cc_10 N_NET27_13 N_A1_9 0.000814008f
cc_11 N_NET27_1 N_MM0_g 0.0010065f
cc_12 N_NET27_10 N_MM0_g 0.0340907f
cc_13 N_NET27_16 N_A2_6 0.000459185f
cc_14 N_NET27_10 N_A2_1 0.000649858f
cc_15 N_NET27_1 N_A2_4 0.000818807f
cc_16 N_NET27_1 N_MM10_g 0.00139113f
cc_17 N_NET27_13 N_A2_6 0.0043587f
cc_18 N_NET27_10 N_MM10_g 0.0342403f
cc_19 N_NET27_16 N_A3_4 0.000555301f
cc_20 N_NET27_11 N_A3_1 0.000677097f
cc_21 N_NET27_2 N_MM13_g 0.000853166f
cc_22 N_NET27_2 N_A3_4 0.00106619f
cc_23 N_NET27_11 N_MM13_g 0.0342383f
cc_24 N_NET27_11 N_B2_1 0.000773397f
cc_25 N_NET27_2 N_MM11_g 0.00085062f
cc_26 N_NET27_15 N_B2_4 0.00102753f
cc_27 N_NET27_2 N_B2_4 0.00125228f
cc_28 N_NET27_11 N_MM11_g 0.0337722f
cc_29 N_NET27_12 N_B1_1 0.000838278f
cc_30 N_NET27_3 N_MM8_g 0.00118443f
cc_31 N_NET27_15 N_B1_6 0.00448457f
cc_32 N_NET27_12 N_MM8_g 0.034618f
x_PM_AO322x2_ASAP7_75t_R%A3 VSS A3 N_MM13_g N_A3_1 N_A3_4
+ PM_AO322x2_ASAP7_75t_R%A3
cc_33 N_MM13_g N_A2_1 0.00089395f
cc_34 N_A3_1 N_A2_1 0.00125981f
cc_35 N_A3_4 N_A2_4 0.00382115f
cc_36 N_MM13_g N_MM10_g 0.00571941f
x_PM_AO322x2_ASAP7_75t_R%B2 VSS B2 N_MM11_g N_B2_1 N_B2_4
+ PM_AO322x2_ASAP7_75t_R%B2
cc_37 N_B2_1 N_MM13_g 0.000840302f
cc_38 N_B2_4 N_A3_4 0.0031714f
cc_39 N_MM11_g N_MM13_g 0.0040401f
x_PM_AO322x2_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_AO322x2_ASAP7_75t_R%noxref_18
cc_40 N_noxref_18_1 N_MM0_g 0.00215469f
cc_41 N_noxref_18_1 N_NET25_4 0.000512917f
cc_42 N_noxref_18_1 N_NET25_21 0.0367316f
x_PM_AO322x2_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_AO322x2_ASAP7_75t_R%noxref_19
cc_43 N_noxref_19_1 N_MM0_g 0.00223056f
cc_44 N_noxref_19_1 N_NET25_21 0.00050014f
cc_45 N_noxref_19_1 N_noxref_18_1 0.00176268f
x_PM_AO322x2_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_AO322x2_ASAP7_75t_R%noxref_20
cc_46 N_noxref_20_1 N_MM8_g 0.00348568f
cc_47 N_noxref_20_1 N_NET25_6 0.000107789f
cc_48 N_noxref_20_1 N_NET25_27 0.000132998f
cc_49 N_noxref_20_1 N_NET25_5 0.00046063f
cc_50 N_noxref_20_1 N_NET25_22 0.027357f
cc_51 N_noxref_20_1 N_NET27_12 0.000493777f
x_PM_AO322x2_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_AO322x2_ASAP7_75t_R%noxref_22
cc_52 N_noxref_22_1 N_MM9_g 0.00337006f
cc_53 N_noxref_22_1 N_NET25_22 6.30831e-20
cc_54 N_noxref_22_1 N_NET25_7 6.35298e-20
cc_55 N_noxref_22_1 N_NET25_24 9.53519e-20
cc_56 N_noxref_22_1 N_NET25_5 0.000121355f
cc_57 N_noxref_22_1 N_NET25_27 0.000170967f
cc_58 N_noxref_22_1 N_NET25_6 0.000435954f
cc_59 N_noxref_22_1 N_NET25_23 0.0275503f
cc_60 N_noxref_22_1 N_noxref_20_1 0.00777269f
cc_61 N_noxref_22_1 N_noxref_21_1 0.000474205f
x_PM_AO322x2_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_AO322x2_ASAP7_75t_R%noxref_23
cc_62 N_noxref_23_1 N_MM9_g 0.0015021f
cc_63 N_noxref_23_1 N_NET25_7 0.000412142f
cc_64 N_noxref_23_1 N_NET25_24 0.0370655f
cc_65 N_noxref_23_1 N_NET27_12 0.000558572f
cc_66 N_noxref_23_1 N_noxref_20_1 0.000475053f
cc_67 N_noxref_23_1 N_noxref_21_1 0.00766461f
cc_68 N_noxref_23_1 N_noxref_22_1 0.00135518f
x_PM_AO322x2_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_AO322x2_ASAP7_75t_R%noxref_24
cc_69 N_noxref_24_1 N_MM12_g 0.00345649f
cc_70 N_noxref_24_1 N_NET25_8 6.35008e-20
cc_71 N_noxref_24_1 N_NET25_30 8.32922e-20
cc_72 N_noxref_24_1 N_NET25_25 0.000753921f
cc_73 N_noxref_24_1 N_Y_13 0.000719164f
x_PM_AO322x2_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_AO322x2_ASAP7_75t_R%noxref_21
cc_74 N_noxref_21_1 N_MM8_g 0.00155529f
cc_75 N_noxref_21_1 N_NET25_7 0.000128969f
cc_76 N_noxref_21_1 N_NET25_24 0.000724793f
cc_77 N_noxref_21_1 N_NET27_12 0.0355971f
cc_78 N_noxref_21_1 N_noxref_20_1 0.00135647f
x_PM_AO322x2_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_AO322x2_ASAP7_75t_R%noxref_25
cc_79 N_noxref_25_1 N_MM12_g 0.0014939f
cc_80 N_noxref_25_1 N_NET25_30 6.1926e-20
cc_81 N_noxref_25_1 N_NET25_8 0.000417759f
cc_82 N_noxref_25_1 N_NET25_25 0.0370169f
cc_83 N_noxref_25_1 N_Y_15 0.000680212f
cc_84 N_noxref_25_1 N_noxref_24_1 0.00134382f
x_PM_AO322x2_ASAP7_75t_R%C1 VSS C1 N_MM9_g N_C1_1 N_C1_4
+ PM_AO322x2_ASAP7_75t_R%C1
x_PM_AO322x2_ASAP7_75t_R%noxref_26 VSS N_noxref_26_1
+ PM_AO322x2_ASAP7_75t_R%noxref_26
cc_85 N_noxref_26_1 N_MM17_g 0.00168443f
cc_86 N_noxref_26_1 N_Y_13 0.0372267f
cc_87 N_noxref_26_1 N_noxref_24_1 0.00771487f
x_PM_AO322x2_ASAP7_75t_R%A2 VSS A2 N_MM10_g N_A2_6 N_A2_5 N_A2_1 N_A2_4
+ PM_AO322x2_ASAP7_75t_R%A2
cc_88 N_A2_6 N_A1_6 0.000508593f
cc_89 N_A2_5 N_A1_6 0.000524001f
cc_90 N_A2_1 N_A1_1 0.00199146f
cc_91 N_A2_4 N_A1_6 0.00267807f
cc_92 N_MM10_g N_MM0_g 0.00637371f
x_PM_AO322x2_ASAP7_75t_R%C2 VSS C2 N_MM12_g N_C2_1 N_C2_4 N_C2_5
+ PM_AO322x2_ASAP7_75t_R%C2
cc_93 N_C2_1 N_C1_1 0.0021889f
cc_94 N_C2_4 N_C1_4 0.00339117f
cc_95 N_MM12_g N_MM9_g 0.00714369f
x_PM_AO322x2_ASAP7_75t_R%A1 VSS A1 N_MM0_g N_A1_6 N_A1_1 N_A1_4 N_A1_7 N_A1_9
+ PM_AO322x2_ASAP7_75t_R%A1
x_PM_AO322x2_ASAP7_75t_R%noxref_27 VSS N_noxref_27_1
+ PM_AO322x2_ASAP7_75t_R%noxref_27
cc_96 N_noxref_27_1 N_NET25_30 7.46358e-20
cc_97 N_noxref_27_1 N_NET25_25 8.81178e-20
cc_98 N_noxref_27_1 N_NET25_8 0.000133874f
cc_99 N_noxref_27_1 N_MM17_g 0.00193225f
cc_100 N_noxref_27_1 N_Y_15 0.0372381f
cc_101 N_noxref_27_1 N_noxref_24_1 0.000469705f
cc_102 N_noxref_27_1 N_noxref_25_1 0.00766894f
cc_103 N_noxref_27_1 N_noxref_26_1 0.00123745f
x_PM_AO322x2_ASAP7_75t_R%noxref_29 VSS N_noxref_29_1
+ PM_AO322x2_ASAP7_75t_R%noxref_29
cc_104 N_noxref_29_1 N_MM17@2_g 0.00149728f
cc_105 N_noxref_29_1 N_Y_16 0.0380229f
cc_106 N_noxref_29_1 N_noxref_28_1 0.0017637f
x_PM_AO322x2_ASAP7_75t_R%B1 VSS B1 N_MM8_g N_B1_1 N_B1_4 N_B1_5 N_B1_6
+ PM_AO322x2_ASAP7_75t_R%B1
cc_107 N_B1_1 N_B2_1 0.00206347f
cc_108 N_B1_4 N_B2_4 0.00294395f
cc_109 N_MM8_g N_MM11_g 0.00735533f
x_PM_AO322x2_ASAP7_75t_R%noxref_28 VSS N_noxref_28_1
+ PM_AO322x2_ASAP7_75t_R%noxref_28
cc_110 N_noxref_28_1 N_MM17@2_g 0.00149242f
cc_111 N_noxref_28_1 N_Y_14 0.0382827f
x_PM_AO322x2_ASAP7_75t_R%NET53 VSS N_MM11_d N_MM8_d N_MM9_s N_MM12_s N_NET53_7
+ N_NET53_1 N_NET53_8 N_NET53_2 N_NET53_9 PM_AO322x2_ASAP7_75t_R%NET53
cc_112 N_NET53_7 N_B2_1 0.000736705f
cc_113 N_NET53_1 N_MM11_g 0.000900896f
cc_114 N_NET53_7 N_MM11_g 0.0336648f
cc_115 N_NET53_7 N_B1_1 0.000657217f
cc_116 N_NET53_1 N_MM8_g 0.000948374f
cc_117 N_NET53_7 N_MM8_g 0.0340088f
cc_118 N_NET53_8 N_C1_1 0.000629309f
cc_119 N_NET53_2 N_MM9_g 0.000903421f
cc_120 N_NET53_8 N_MM9_g 0.0335877f
cc_121 N_NET53_8 N_C2_1 0.000612877f
cc_122 N_NET53_2 N_MM12_g 0.000903447f
cc_123 N_NET53_8 N_MM12_g 0.0335515f
cc_124 N_NET53_9 N_NET25_25 0.00064924f
cc_125 N_NET53_9 N_NET25_8 0.000229556f
cc_126 N_NET53_9 N_NET25_27 0.000358688f
cc_127 N_NET53_8 N_NET25_24 0.00058837f
cc_128 N_NET53_2 N_NET25_28 0.000709666f
cc_129 N_NET53_9 N_NET25_7 0.000709893f
cc_130 N_NET53_8 N_NET25_25 0.00112295f
cc_131 N_NET53_2 N_NET25_7 0.00166751f
cc_132 N_NET53_9 N_NET25_28 0.00400784f
cc_133 N_NET53_2 N_NET25_8 0.00434339f
cc_134 N_NET53_9 N_NET25_32 0.00646949f
cc_135 N_NET53_7 N_NET27_12 0.00170468f
cc_136 N_NET53_1 N_NET27_15 0.000798854f
cc_137 N_NET53_1 N_NET27_2 0.00124098f
cc_138 N_NET53_1 N_NET27_3 0.00472851f
cc_139 N_NET53_9 N_NET27_15 0.00982371f
x_PM_AO322x2_ASAP7_75t_R%Y VSS Y N_MM16_d N_MM16@2_d N_MM17@2_d N_MM17_d N_Y_14
+ N_Y_18 N_Y_2 N_Y_16 N_Y_13 N_Y_15 N_Y_1 N_Y_17 N_Y_3 N_Y_4 N_Y_19
+ PM_AO322x2_ASAP7_75t_R%Y
cc_140 N_Y_14 N_NET25_8 0.000284216f
cc_141 N_Y_14 N_NET25_25 8.17071e-20
cc_142 N_Y_14 N_NET25_28 0.000114553f
cc_143 N_Y_14 N_NET25_33 0.000134001f
cc_144 N_Y_14 N_MM17_g 0.000351838f
cc_145 N_Y_18 N_NET25_34 0.00029382f
cc_146 N_Y_2 N_NET25_29 0.000311808f
cc_147 N_Y_16 N_MM17@2_g 0.0154881f
cc_148 N_Y_13 N_MM17_g 0.053766f
cc_149 N_Y_15 N_MM17_g 0.0157366f
cc_150 N_Y_1 N_NET25_1 0.000713963f
cc_151 N_Y_17 N_NET25_30 0.000905524f
cc_152 N_Y_3 N_MM17@2_g 0.00110283f
cc_153 N_Y_4 N_MM17@2_g 0.00111187f
cc_154 N_Y_3 N_NET25_1 0.00112191f
cc_155 N_Y_18 N_NET25_30 0.00115441f
cc_156 N_Y_1 N_MM17_g 0.00158334f
cc_157 N_Y_2 N_MM17_g 0.00187326f
cc_158 N_Y_19 N_NET25_30 0.00189932f
cc_159 N_Y_16 N_NET25_1 0.00338723f
cc_160 N_Y_1 N_NET25_30 0.0042577f
cc_161 N_Y_14 N_MM17@2_g 0.0540443f
x_PM_AO322x2_ASAP7_75t_R%NET25 VSS N_MM17_g N_MM17@2_g N_MM12_d N_MM9_d N_MM5_d
+ N_MM3_d N_MM0_d N_NET25_4 N_NET25_21 N_NET25_26 N_NET25_5 N_NET25_22
+ N_NET25_32 N_NET25_27 N_NET25_7 N_NET25_6 N_NET25_23 N_NET25_31 N_NET25_28
+ N_NET25_24 N_NET25_8 N_NET25_30 N_NET25_33 N_NET25_29 N_NET25_25 N_NET25_34
+ N_NET25_1 PM_AO322x2_ASAP7_75t_R%NET25
cc_162 N_NET25_4 N_MM0_g 0.00356744f
cc_163 N_NET25_4 N_A1_4 0.000558482f
cc_164 N_NET25_21 N_A1_1 0.0010153f
cc_165 N_NET25_26 N_A1_6 0.00156624f
cc_166 N_NET25_26 N_A1_7 0.00203399f
cc_167 N_NET25_21 N_MM0_g 0.0356261f
cc_168 N_NET25_21 N_A2_5 0.000623558f
cc_169 N_NET25_4 N_A2_5 0.000409627f
cc_170 N_NET25_26 N_A2_4 0.000436508f
cc_171 N_NET25_26 N_A2_5 0.00533276f
cc_172 N_NET25_21 N_A3_4 8.07144e-20
cc_173 N_NET25_26 N_A3_4 0.00270099f
cc_174 N_NET25_5 N_B2_4 0.000166659f
cc_175 N_NET25_22 N_B2_4 0.000226943f
cc_176 N_NET25_26 N_B2_4 0.00281121f
cc_177 N_NET25_5 N_MM8_g 0.00148463f
cc_178 N_NET25_32 N_MM8_g 8.44559e-20
cc_179 N_NET25_5 N_B1_5 0.00033577f
cc_180 N_NET25_27 N_B1_6 0.000340334f
cc_181 N_NET25_22 N_B1_1 0.000400828f
cc_182 N_NET25_27 N_B1_5 0.000811224f
cc_183 N_NET25_5 N_B1_4 0.000879717f
cc_184 N_NET25_26 N_B1_5 0.00538112f
cc_185 N_NET25_22 N_MM8_g 0.0256076f
cc_186 N_NET25_32 N_MM9_g 5.7388e-20
cc_187 N_NET25_7 N_MM9_g 0.00120211f
cc_188 N_NET25_6 N_MM9_g 0.00117101f
cc_189 N_NET25_23 N_MM9_g 0.0113269f
cc_190 N_NET25_31 N_C1_4 0.000509061f
cc_191 N_NET25_7 N_C1_1 0.000810763f
cc_192 N_NET25_28 N_C1_4 0.00115664f
cc_193 N_NET25_24 N_C1_1 0.00128478f
cc_194 N_NET25_27 N_C1_4 0.00620254f
cc_195 N_NET25_24 N_MM9_g 0.0491325f
cc_196 N_NET25_6 N_MM12_g 0.000281056f
cc_197 N_NET25_23 N_MM12_g 8.4492e-20
cc_198 N_NET25_31 N_MM12_g 0.000112336f
cc_199 N_NET25_8 N_MM12_g 0.00118906f
cc_200 N_NET25_27 N_MM12_g 0.000149679f
cc_201 N_NET25_30 N_C2_5 0.00045582f
cc_202 N_NET25_33 N_C2_5 0.000576363f
cc_203 N_NET25_8 N_C2_1 0.000647397f
cc_204 N_NET25_29 N_C2_4 0.000677347f
cc_205 N_NET25_25 N_C2_1 0.000968643f
cc_206 N_NET25_28 N_C2_4 0.00116098f
cc_207 N_NET25_33 N_C2_4 0.00342002f
cc_208 N_NET25_25 N_MM12_g 0.0354021f
*END of AO322x2_ASAP7_75t_R.pxi
.ENDS
** Design:	AO32x1_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AO32x1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AO32x1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AO32x1_ASAP7_75t_R%NET26 VSS 2 3 1
c1 1 VSS 0.000886139f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0540 $X2=0.3240 $Y2=0.0540
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0540 $X2=0.3240 $Y2=0.0540
.ends

.subckt PM_AO32x1_ASAP7_75t_R%NET24 VSS 2 3 1
c1 1 VSS 0.000933094f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2160 $Y2=0.0675
.ends

.subckt PM_AO32x1_ASAP7_75t_R%NET25 VSS 2 3 1
c1 1 VSS 0.000882053f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_AO32x1_ASAP7_75t_R%A3 VSS 8 3 4 1
c1 1 VSS 0.00657711f
c2 3 VSS 0.0833873f
c3 4 VSS 0.00566034f
r1 8 7 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1755 $X2=0.1350 $Y2=0.1595
r2 4 7 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1595
r3 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r4 1 4 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AO32x1_ASAP7_75t_R%A1 VSS 9 3 1 4
c1 1 VSS 0.00509049f
c2 3 VSS 0.0347438f
c3 4 VSS 0.00419664f
r1 9 8 1.51573 $w=1.3e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1765 $X2=0.2430 $Y2=0.1700
r2 7 8 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1540 $X2=0.2430 $Y2=0.1700
r3 6 7 4.4306 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1540
r4 4 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0980 $X2=0.2430 $Y2=0.1350
r5 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r6 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AO32x1_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00491342f
.ends

.subckt PM_AO32x1_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00475628f
.ends

.subckt PM_AO32x1_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.0319497f
.ends

.subckt PM_AO32x1_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.00523981f
.ends

.subckt PM_AO32x1_ASAP7_75t_R%A2 VSS 6 3 4 1
c1 1 VSS 0.00442823f
c2 3 VSS 0.0353019f
c3 4 VSS 0.00385394f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.0980
r2 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AO32x1_ASAP7_75t_R%Y VSS 21 14 29 7 2 1 8 12 9
c1 1 VSS 0.00745924f
c2 2 VSS 0.00861946f
c3 7 VSS 0.00373059f
c4 8 VSS 0.00370175f
c5 9 VSS 0.00290117f
c6 10 VSS 0.00102018f
c7 11 VSS 0.00606192f
c8 12 VSS 0.0031465f
r1 29 28 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r2 8 28 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r3 2 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0535 $Y2=0.2340
r4 24 25 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.2340 $X2=0.0535 $Y2=0.2340
r5 11 23 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0270 $Y2=0.2125
r6 11 24 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0405 $Y2=0.2340
r7 22 23 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1880 $X2=0.0270 $Y2=0.2125
r8 21 22 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1755 $X2=0.0270 $Y2=0.1880
r9 21 20 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1755 $X2=0.0270 $Y2=0.1595
r10 19 20 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1350 $X2=0.0270 $Y2=0.1595
r11 9 18 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1035 $X2=0.0270 $Y2=0.0720
r12 9 19 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1035 $X2=0.0270 $Y2=0.1350
r13 10 17 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0405 $Y=0.0720 $X2=0.0540 $Y2=0.0720
r14 10 18 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0405 $Y=0.0720 $X2=0.0270 $Y2=0.0720
r15 16 17 1.50137 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0540 $Y=0.0605 $X2=0.0540 $Y2=0.0720
r16 15 16 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.0490 $X2=0.0540 $Y2=0.0605
r17 12 15 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.0370 $X2=0.0540 $Y2=0.0490
r18 1 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0540 $Y2=0.0490
r19 14 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r20 7 13 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r21 2 8 1e-05
r22 1 7 1e-05
.ends

.subckt PM_AO32x1_ASAP7_75t_R%B1 VSS 6 3 1 4
c1 1 VSS 0.00510527f
c2 3 VSS 0.00797436f
c3 4 VSS 0.00344301f
r1 7 8 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1230 $X2=0.2970 $Y2=0.1350
r2 6 7 0.816164 $w=1.3e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1195 $X2=0.2970 $Y2=0.1230
r3 6 4 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1195 $X2=0.2970 $Y2=0.0945
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_AO32x1_ASAP7_75t_R%B2 VSS 6 3 1 4
c1 1 VSS 0.00438202f
c2 3 VSS 0.0345997f
c3 4 VSS 0.00337044f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.0980
r2 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
.ends

.subckt PM_AO32x1_ASAP7_75t_R%NET10 VSS 15 18 34 35 37 13 12 3 2 1 10 11
c1 1 VSS 0.0088652f
c2 2 VSS 0.00610029f
c3 3 VSS 0.00531872f
c4 10 VSS 0.00397424f
c5 11 VSS 0.00290976f
c6 12 VSS 0.00234167f
c7 13 VSS 0.0218907f
r1 12 3 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2160 $X2=0.3760 $Y2=0.2160
r2 37 12 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2160 $X2=0.3635 $Y2=0.2160
r3 35 33 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2160 $X2=0.1765 $Y2=0.2160
r4 1 33 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2160 $X2=0.1765 $Y2=0.2160
r5 10 1 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1620 $Y2=0.2160
r6 34 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r7 3 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2160
+ $X2=0.3780 $Y2=0.2340
r8 1 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r9 29 30 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3395
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r10 28 29 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3080
+ $Y=0.2340 $X2=0.3395 $Y2=0.2340
r11 27 28 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.2340 $X2=0.3080 $Y2=0.2340
r12 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r13 23 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r14 22 23 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.1890 $Y2=0.2340
r15 21 22 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r16 20 27 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2835
+ $Y=0.2340 $X2=0.2970 $Y2=0.2340
r17 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.2835 $Y2=0.2340
r18 13 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r19 13 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.2340 $X2=0.2430 $Y2=0.2340
r20 2 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2160
+ $X2=0.2700 $Y2=0.2340
r21 18 17 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2160 $X2=0.2845 $Y2=0.2160
r22 16 17 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2800 $Y=0.2160 $X2=0.2845 $Y2=0.2160
r23 2 16 0.222222 $w=5.4e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2680 $Y=0.2160 $X2=0.2800 $Y2=0.2160
r24 11 2 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2160 $X2=0.2680 $Y2=0.2160
r25 15 11 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2160 $X2=0.2555 $Y2=0.2160
.ends

.subckt PM_AO32x1_ASAP7_75t_R%NET08 VSS 9 53 54 68 69 1 15 14 18 3 11 10 4 13
+ 16 17 19 21
c1 1 VSS 0.00352702f
c2 3 VSS 0.00540662f
c3 4 VSS 0.00295827f
c4 9 VSS 0.0803153f
c5 10 VSS 0.0027828f
c6 11 VSS 0.000882853f
c7 12 VSS 0.000219052f
c8 13 VSS 0.0030055f
c9 14 VSS 0.00241795f
c10 15 VSS 0.0281216f
c11 16 VSS 0.00108843f
c12 17 VSS 0.00545647f
c13 18 VSS 0.000837929f
c14 19 VSS 0.00320117f
c15 20 VSS 0.003734f
c16 21 VSS 0.00119859f
r1 69 67 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2160 $X2=0.3385 $Y2=0.2160
r2 4 67 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2160 $X2=0.3385 $Y2=0.2160
r3 13 4 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2160 $X2=0.3240 $Y2=0.2160
r4 68 13 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2160 $X2=0.3095 $Y2=0.2160
r5 4 64 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2160
+ $X2=0.3240 $Y2=0.1980
r6 64 65 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1980 $X2=0.3375 $Y2=0.1980
r7 62 65 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1980 $X2=0.3375 $Y2=0.1980
r8 61 62 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3760
+ $Y=0.1980 $X2=0.3510 $Y2=0.1980
r9 16 21 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3940 $Y=0.1980 $X2=0.4050 $Y2=0.1980
r10 16 61 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3940
+ $Y=0.1980 $X2=0.3760 $Y2=0.1980
r11 21 60 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.1980 $X2=0.4050 $Y2=0.1765
r12 59 60 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1170 $X2=0.4050 $Y2=0.1765
r13 17 20 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.0575 $X2=0.4050 $Y2=0.0360
r14 17 59 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0575 $X2=0.4050 $Y2=0.1170
r15 57 58 0.264706 $w=1.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2800 $Y=0.0725 $X2=0.2845 $Y2=0.0725
r16 3 57 0.705882 $w=1.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2680 $Y=0.0725 $X2=0.2800 $Y2=0.0725
r17 12 3 0.735294 $w=1.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0725 $X2=0.2680 $Y2=0.0725
r18 11 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0945 $X2=0.2680 $Y2=0.0945
r19 54 52 0.0675676 $w=3.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0455 $X2=0.2845 $Y2=0.0455
r20 3 52 0.391892 $w=3.7e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.0455 $X2=0.2845 $Y2=0.0455
r21 3 58 0.471383 $w=3.35517e-08 $l=3.06472e-08 $layer=N_src_drn
+ $thickness=1e-09 $X=0.2700 $Y=0.0455 $X2=0.2845 $Y2=0.0725
r22 10 3 0.391892 $w=3.7e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0455 $X2=0.2700 $Y2=0.0455
r23 53 10 0.0675676 $w=3.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0455 $X2=0.2555 $Y2=0.0455
r24 20 49 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.0360 $X2=0.3780 $Y2=0.0360
r25 3 43 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0540
+ $X2=0.2700 $Y2=0.0360
r26 48 49 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r27 47 48 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3260
+ $Y=0.0360 $X2=0.3510 $Y2=0.0360
r28 46 47 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3080
+ $Y=0.0360 $X2=0.3260 $Y2=0.0360
r29 45 46 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.3080 $Y2=0.0360
r30 44 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2835
+ $Y=0.0360 $X2=0.2970 $Y2=0.0360
r31 43 44 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.2835 $Y2=0.0360
r32 42 43 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r33 41 42 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2565 $Y2=0.0360
r34 40 41 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r35 39 40 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r36 38 39 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1640
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r37 37 38 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1460
+ $Y=0.0360 $X2=0.1640 $Y2=0.0360
r38 36 37 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1460 $Y2=0.0360
r39 15 19 2.65995 $w=1.48966e-08 $l=1.83371e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1170 $Y=0.0360 $X2=0.0990 $Y2=0.0395
r40 15 36 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1170
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r41 19 34 3.47612 $w=1.45278e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0990 $Y=0.0395 $X2=0.0990 $Y2=0.0575
r42 33 34 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0990
+ $Y=0.0755 $X2=0.0990 $Y2=0.0575
r43 14 32 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0990 $Y=0.1035 $X2=0.0990 $Y2=0.1350
r44 14 33 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0990
+ $Y=0.1035 $X2=0.0990 $Y2=0.0755
r45 31 32 1.50137 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0875 $Y=0.1350 $X2=0.0990 $Y2=0.1350
r46 30 31 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0765
+ $Y=0.1350 $X2=0.0875 $Y2=0.1350
r47 28 30 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0675
+ $Y=0.1350 $X2=0.0765 $Y2=0.1350
r48 18 28 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0650
+ $Y=0.1350 $X2=0.0675 $Y2=0.1350
r49 23 27 1.07884 $w=2.10429e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0880 $Y=0.1350 $X2=0.0915 $Y2=0.1350
r50 1 23 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.0780
+ $Y=0.1350 $X2=0.0880 $Y2=0.1350
r51 9 1 2.14279 $w=1.42588e-07 $l=3e-09 $layer=LIG $thickness=5.27059e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0780 $Y2=0.1350
r52 1 25 3.00957 $w=2.05111e-08 $l=9e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0780 $Y=0.1350 $X2=0.0690 $Y2=0.1350
r53 1 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0780 $Y=0.1350
+ $X2=0.0765 $Y2=0.1350
r54 9 25 1.49611 $w=1.91717e-07 $l=1.2e-08 $layer=LIG $thickness=5.46667e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0690 $Y2=0.1350
r55 9 27 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.0810 $Y=0.1350 $X2=0.0915 $Y2=0.1350
.ends


*
.SUBCKT AO32x1_ASAP7_75t_R VSS VDD A3 A2 A1 B1 B2 Y
*
* VSS VSS
* VDD VDD
* A3 A3
* A2 A2
* A1 A1
* B1 B1
* B2 B2
* Y Y
*
*

MM21 N_MM21_d N_MM21_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM0_g N_MM0_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM13 N_MM13_d N_MM14_g N_MM13_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM18 N_MM18_d N_MM15_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM20 N_MM20_d N_MM21_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1 N_MM1_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM14 N_MM14_d N_MM14_g N_MM14_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM15 N_MM15_d N_MM15_g N_MM15_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2


*include "AO32x1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AO32x1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AO32x1_ASAP7_75t_R%NET26 VSS N_MM13_s N_MM18_d N_NET26_1
+ PM_AO32x1_ASAP7_75t_R%NET26
cc_1 N_NET26_1 N_MM14_g 0.0125205f
cc_2 N_NET26_1 N_MM15_g 0.0125767f
x_PM_AO32x1_ASAP7_75t_R%NET24 VSS N_MM2_d N_MM0_s N_NET24_1
+ PM_AO32x1_ASAP7_75t_R%NET24
cc_3 N_NET24_1 N_MM2_g 0.0173727f
cc_4 N_NET24_1 N_MM0_g 0.0173742f
x_PM_AO32x1_ASAP7_75t_R%NET25 VSS N_MM3_d N_MM2_s N_NET25_1
+ PM_AO32x1_ASAP7_75t_R%NET25
cc_5 N_NET25_1 N_MM3_g 0.017285f
cc_6 N_NET25_1 N_MM2_g 0.017415f
x_PM_AO32x1_ASAP7_75t_R%A3 VSS A3 N_MM3_g N_A3_4 N_A3_1 PM_AO32x1_ASAP7_75t_R%A3
cc_7 N_A3_4 N_NET08_1 0.00102123f
cc_8 N_A3_4 N_NET08_15 0.00106307f
cc_9 N_A3_4 N_NET08_14 0.00238946f
cc_10 N_MM3_g N_MM21_g 0.00337282f
cc_11 N_A3_4 N_NET08_18 0.00593514f
x_PM_AO32x1_ASAP7_75t_R%A1 VSS A1 N_MM0_g N_A1_1 N_A1_4 PM_AO32x1_ASAP7_75t_R%A1
cc_12 N_MM0_g N_NET08_10 0.0101496f
cc_13 N_MM0_g N_NET08_3 0.00184263f
cc_14 N_A1_1 N_NET08_10 0.000852878f
cc_15 N_A1_4 N_NET08_15 0.00133436f
cc_16 N_A1_4 N_NET08_3 0.00220822f
cc_17 N_MM0_g N_NET08_11 0.0253505f
cc_18 N_A1_1 N_A2_1 0.00158991f
cc_19 N_A1_4 N_A2_4 0.00489005f
cc_20 N_MM0_g N_MM2_g 0.00822947f
x_PM_AO32x1_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_AO32x1_ASAP7_75t_R%noxref_14
cc_21 N_noxref_14_1 N_MM21_g 0.00147708f
cc_22 N_noxref_14_1 N_Y_7 0.0382977f
x_PM_AO32x1_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_AO32x1_ASAP7_75t_R%noxref_15
cc_23 N_noxref_15_1 N_MM21_g 0.00147108f
cc_24 N_noxref_15_1 N_Y_8 0.0384779f
cc_25 N_noxref_15_1 N_noxref_14_1 0.00177376f
x_PM_AO32x1_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_AO32x1_ASAP7_75t_R%noxref_16
cc_26 N_noxref_16_1 N_NET08_17 0.000941907f
cc_27 N_noxref_16_1 N_MM15_g 0.00369472f
x_PM_AO32x1_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_AO32x1_ASAP7_75t_R%noxref_17
cc_28 N_noxref_17_1 N_NET08_13 0.000921903f
cc_29 N_noxref_17_1 N_MM15_g 0.00366778f
cc_30 N_noxref_17_1 N_NET10_12 0.026675f
cc_31 N_noxref_17_1 N_noxref_16_1 0.00205591f
x_PM_AO32x1_ASAP7_75t_R%A2 VSS A2 N_MM2_g N_A2_4 N_A2_1 PM_AO32x1_ASAP7_75t_R%A2
cc_32 N_A2_4 N_NET08_3 0.000277359f
cc_33 N_MM2_g N_NET08_11 0.000445271f
cc_34 N_A2_4 N_NET08_15 0.00147255f
cc_35 N_A2_4 N_NET08_18 0.002083f
cc_36 N_A2_1 N_A3_1 0.00167206f
cc_37 N_A2_4 N_A3_4 0.00502869f
cc_38 N_MM2_g N_MM3_g 0.00831349f
x_PM_AO32x1_ASAP7_75t_R%Y VSS Y N_MM21_d N_MM20_d N_Y_7 N_Y_2 N_Y_1 N_Y_8
+ N_Y_12 N_Y_9 PM_AO32x1_ASAP7_75t_R%Y
cc_39 N_Y_7 N_NET08_14 0.000359658f
cc_40 N_Y_7 N_NET08_19 0.000520237f
cc_41 N_Y_2 N_NET08_1 0.00105873f
cc_42 N_Y_2 N_MM21_g 0.00119804f
cc_43 N_Y_1 N_MM21_g 0.0013932f
cc_44 N_Y_8 N_NET08_1 0.00207105f
cc_45 N_Y_12 N_NET08_14 0.00320523f
cc_46 N_Y_9 N_NET08_18 0.00342571f
cc_47 N_Y_8 N_MM21_g 0.0153061f
cc_48 N_Y_7 N_MM21_g 0.0547699f
x_PM_AO32x1_ASAP7_75t_R%B1 VSS B1 N_MM14_g N_B1_1 N_B1_4
+ PM_AO32x1_ASAP7_75t_R%B1
cc_49 N_MM14_g N_NET08_4 0.000679542f
cc_50 N_MM14_g N_NET08_11 0.00561202f
cc_51 N_MM14_g N_NET08_13 0.0112202f
cc_52 N_B1_1 N_NET08_3 0.000439559f
cc_53 N_B1_4 N_NET08_16 0.000584307f
cc_54 N_B1_1 N_NET08_10 0.00108766f
cc_55 N_B1_4 N_NET08_15 0.00130651f
cc_56 N_MM14_g N_NET08_3 0.00156557f
cc_57 N_B1_4 N_NET08_3 0.00256701f
cc_58 N_MM14_g N_NET08_10 0.0442556f
cc_59 N_B1_1 N_A1_1 0.00119468f
cc_60 N_B1_4 N_A1_4 0.00372299f
cc_61 N_MM14_g N_MM0_g 0.00623914f
x_PM_AO32x1_ASAP7_75t_R%B2 VSS B2 N_MM15_g N_B2_1 N_B2_4
+ PM_AO32x1_ASAP7_75t_R%B2
cc_62 N_MM15_g N_NET08_3 0.000261031f
cc_63 N_MM15_g N_NET08_4 0.000409849f
cc_64 N_B2_1 N_NET08_17 0.000620124f
cc_65 N_B2_1 N_NET08_13 0.000679825f
cc_66 N_B2_4 N_NET08_16 0.00118939f
cc_67 N_B2_4 N_NET08_15 0.00125089f
cc_68 N_B2_4 N_NET08_17 0.00651582f
cc_69 N_MM15_g N_NET08_13 0.0258904f
cc_70 N_B2_1 N_B1_1 0.00160947f
cc_71 N_B2_4 N_B1_4 0.00351132f
cc_72 N_MM15_g N_MM14_g 0.00966855f
x_PM_AO32x1_ASAP7_75t_R%NET10 VSS N_MM5_d N_MM14_s N_MM4_d N_MM1_d N_MM15_s
+ N_NET10_13 N_NET10_12 N_NET10_3 N_NET10_2 N_NET10_1 N_NET10_10 N_NET10_11
+ PM_AO32x1_ASAP7_75t_R%NET10
cc_73 N_NET10_13 N_NET08_13 0.000424985f
cc_74 N_NET10_13 N_NET08_17 0.000469233f
cc_75 N_NET10_12 N_NET08_13 0.00135023f
cc_76 N_NET10_3 N_NET08_16 0.000567048f
cc_77 N_NET10_13 N_NET08_21 0.000607077f
cc_78 N_NET10_13 N_NET08_4 0.000741833f
cc_79 N_NET10_2 N_NET08_4 0.00097281f
cc_80 N_NET10_3 N_NET08_4 0.00381824f
cc_81 N_NET10_13 N_NET08_16 0.00869293f
cc_82 N_NET10_1 N_MM3_g 0.000607791f
cc_83 N_NET10_1 N_A3_4 0.000927642f
cc_84 N_NET10_10 N_MM3_g 0.02521f
cc_85 N_NET10_13 N_A2_4 0.00115199f
cc_86 N_NET10_1 N_A2_4 0.00147901f
cc_87 N_NET10_10 N_MM2_g 0.0257083f
cc_88 N_NET10_13 N_A1_4 0.00126809f
cc_89 N_NET10_2 N_A1_4 0.00156282f
cc_90 N_NET10_11 N_MM0_g 0.0255684f
cc_91 N_NET10_2 N_MM14_g 0.000521105f
cc_92 N_NET10_11 N_MM14_g 0.0252458f
cc_93 N_NET10_12 N_MM15_g 0.025642f
x_PM_AO32x1_ASAP7_75t_R%NET08 VSS N_MM21_g N_MM0_d N_MM13_d N_MM14_d N_MM15_d
+ N_NET08_1 N_NET08_15 N_NET08_14 N_NET08_18 N_NET08_3 N_NET08_11 N_NET08_10
+ N_NET08_4 N_NET08_13 N_NET08_16 N_NET08_17 N_NET08_19 N_NET08_21
+ PM_AO32x1_ASAP7_75t_R%NET08
*END of AO32x1_ASAP7_75t_R.pxi
.ENDS
** Design:	AO32x2_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AO32x2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AO32x2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AO32x2_ASAP7_75t_R%NET26 VSS 2 3 1
c1 1 VSS 0.000879847f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0540 $X2=0.3780 $Y2=0.0540
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0540 $X2=0.3780 $Y2=0.0540
.ends

.subckt PM_AO32x2_ASAP7_75t_R%NET24 VSS 2 3 1
c1 1 VSS 0.000931592f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2700 $Y2=0.0675
.ends

.subckt PM_AO32x2_ASAP7_75t_R%NET25 VSS 2 3 1
c1 1 VSS 0.000912507f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2160 $Y2=0.0675
.ends

.subckt PM_AO32x2_ASAP7_75t_R%A3 VSS 8 3 4 1
c1 1 VSS 0.00715445f
c2 3 VSS 0.0835784f
c3 4 VSS 0.00601764f
r1 8 7 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1755 $X2=0.1890 $Y2=0.1595
r2 6 7 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1595
r3 4 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0980 $X2=0.1890 $Y2=0.1350
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r5 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AO32x2_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.0319186f
.ends

.subckt PM_AO32x2_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.00525246f
.ends

.subckt PM_AO32x2_ASAP7_75t_R%A2 VSS 6 3 4 1
c1 1 VSS 0.00452735f
c2 3 VSS 0.0353406f
c3 4 VSS 0.00388481f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.0980
r2 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AO32x2_ASAP7_75t_R%B1 VSS 6 3 1 4
c1 1 VSS 0.00505374f
c2 3 VSS 0.00793429f
c3 4 VSS 0.00335196f
r1 7 8 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1230 $X2=0.3510 $Y2=0.1350
r2 6 7 0.816164 $w=1.3e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1195 $X2=0.3510 $Y2=0.1230
r3 6 4 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1195 $X2=0.3510 $Y2=0.0945
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
.ends

.subckt PM_AO32x2_ASAP7_75t_R%B2 VSS 6 3 1 4
c1 1 VSS 0.00421334f
c2 3 VSS 0.0345361f
c3 4 VSS 0.00332969f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.0980
r2 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
.ends

.subckt PM_AO32x2_ASAP7_75t_R%A1 VSS 10 3 5 1 4
c1 1 VSS 0.00421424f
c2 3 VSS 0.034268f
c3 4 VSS 0.00331497f
c4 5 VSS 0.00260784f
r1 5 11 2.31754 $w=1.6e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1980 $X2=0.2970 $Y2=0.1830
r2 10 11 1.51573 $w=1.3e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1765 $X2=0.2970 $Y2=0.1830
r3 10 9 1.51573 $w=1.3e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1765 $X2=0.2970 $Y2=0.1700
r4 8 9 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1540 $X2=0.2970 $Y2=0.1700
r5 7 8 4.4306 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1540
r6 4 7 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0980 $X2=0.2970 $Y2=0.1350
r7 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r8 1 7 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_AO32x2_ASAP7_75t_R%NET10 VSS 16 17 32 35 37 13 12 3 2 1 10 11
c1 1 VSS 0.00878354f
c2 2 VSS 0.00621102f
c3 3 VSS 0.00531811f
c4 10 VSS 0.00396467f
c5 11 VSS 0.00290933f
c6 12 VSS 0.00234346f
c7 13 VSS 0.021764f
r1 12 3 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2160 $X2=0.4300 $Y2=0.2160
r2 37 12 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2160 $X2=0.4175 $Y2=0.2160
r3 35 34 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2160 $X2=0.3385 $Y2=0.2160
r4 33 34 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3340 $Y=0.2160 $X2=0.3385 $Y2=0.2160
r5 2 33 0.222222 $w=5.4e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3220 $Y=0.2160 $X2=0.3340 $Y2=0.2160
r6 11 2 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2160 $X2=0.3220 $Y2=0.2160
r7 32 11 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2160 $X2=0.3095 $Y2=0.2160
r8 3 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2160
+ $X2=0.4320 $Y2=0.2340
r9 2 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2160
+ $X2=0.3225 $Y2=0.2340
r10 28 29 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3935
+ $Y=0.2340 $X2=0.4320 $Y2=0.2340
r11 27 28 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3620
+ $Y=0.2340 $X2=0.3935 $Y2=0.2340
r12 26 27 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.2340 $X2=0.3620 $Y2=0.2340
r13 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.2340 $X2=0.3510 $Y2=0.2340
r14 24 25 1.39914 $w=1.3e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.3315
+ $Y=0.2340 $X2=0.3375 $Y2=0.2340
r15 23 24 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3225
+ $Y=0.2340 $X2=0.3315 $Y2=0.2340
r16 22 23 4.89699 $w=1.3e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3015
+ $Y=0.2340 $X2=0.3225 $Y2=0.2340
r17 21 22 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.3015 $Y2=0.2340
r18 20 21 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r19 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.2340 $X2=0.2430 $Y2=0.2340
r20 18 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2295 $Y2=0.2340
r21 13 18 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2045
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r22 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2160
+ $X2=0.2160 $Y2=0.2340
r23 16 15 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2160 $X2=0.2305 $Y2=0.2160
r24 1 15 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2160 $X2=0.2305 $Y2=0.2160
r25 10 1 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2160 $X2=0.2160 $Y2=0.2160
r26 17 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2160 $X2=0.2015 $Y2=0.2160
.ends

.subckt PM_AO32x2_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.0424756f
.ends

.subckt PM_AO32x2_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.042393f
.ends

.subckt PM_AO32x2_ASAP7_75t_R%Y VSS 25 17 18 34 35 7 9 8 14 2 1
c1 1 VSS 0.00924144f
c2 2 VSS 0.0107086f
c3 7 VSS 0.00460306f
c4 8 VSS 0.00455725f
c5 9 VSS 0.00580003f
c6 10 VSS 0.00282796f
c7 11 VSS 0.0100495f
c8 12 VSS 0.00154349f
c9 13 VSS 0.00344904f
c10 14 VSS 0.00339879f
r1 35 33 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r2 2 33 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r4 34 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
r5 2 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.2340
r6 29 30 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0960
+ $Y=0.2340 $X2=0.1080 $Y2=0.2340
r7 11 13 7.0955 $w=1.42e-08 $l=3.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.0645
+ $Y=0.2340 $X2=0.0270 $Y2=0.2340
r8 11 29 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0645
+ $Y=0.2340 $X2=0.0960 $Y2=0.2340
r9 13 28 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.2340 $X2=0.0270 $Y2=0.2160
r10 27 28 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.2035 $X2=0.0270 $Y2=0.2160
r11 26 27 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1880 $X2=0.0270 $Y2=0.2035
r12 25 26 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1755 $X2=0.0270 $Y2=0.1880
r13 25 24 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1755 $X2=0.0270 $Y2=0.1595
r14 23 24 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1350 $X2=0.0270 $Y2=0.1595
r15 9 12 5.11339 $w=1.60414e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1060 $X2=0.0270 $Y2=0.0770
r16 9 23 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1060 $X2=0.0270 $Y2=0.1350
r17 12 22 7.0955 $w=1.42e-08 $l=3.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0770 $X2=0.0645 $Y2=0.0770
r18 10 21 1.61797 $w=1.675e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0960 $Y=0.0770 $X2=0.1080 $Y2=0.0770
r19 10 22 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0960
+ $Y=0.0770 $X2=0.0645 $Y2=0.0770
r20 20 21 1.50137 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0655 $X2=0.1080 $Y2=0.0770
r21 19 20 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0540 $X2=0.1080 $Y2=0.0655
r22 14 19 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0410 $X2=0.1080 $Y2=0.0540
r23 1 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1080 $Y2=0.0540
r24 18 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r25 1 16 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r26 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r27 17 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.0935 $Y2=0.0675
.ends

.subckt PM_AO32x2_ASAP7_75t_R%NET08 VSS 9 10 57 58 72 73 1 17 16 21 3 12 11 18
+ 4 14 19 15 20 23
c1 1 VSS 0.00733666f
c2 3 VSS 0.00547294f
c3 4 VSS 0.00281101f
c4 9 VSS 0.0809763f
c5 10 VSS 0.080408f
c6 11 VSS 0.00347027f
c7 12 VSS 0.00159277f
c8 13 VSS 0.000464636f
c9 14 VSS 0.00428404f
c10 15 VSS 0.0017529f
c11 16 VSS 0.00284096f
c12 17 VSS 0.0307894f
c13 18 VSS 0.00160023f
c14 19 VSS 0.00840953f
c15 20 VSS 0.00242296f
c16 21 VSS 0.000356025f
c17 22 VSS 0.00419913f
c18 23 VSS 0.00183073f
r1 73 71 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2160 $X2=0.3925 $Y2=0.2160
r2 4 71 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.2160 $X2=0.3925 $Y2=0.2160
r3 14 4 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2160 $X2=0.3780 $Y2=0.2160
r4 72 14 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2160 $X2=0.3635 $Y2=0.2160
r5 4 68 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2160
+ $X2=0.3780 $Y2=0.1980
r6 68 69 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.1980 $X2=0.3915 $Y2=0.1980
r7 66 69 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1980 $X2=0.3915 $Y2=0.1980
r8 65 66 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4300
+ $Y=0.1980 $X2=0.4050 $Y2=0.1980
r9 18 23 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4480 $Y=0.1980 $X2=0.4590 $Y2=0.1980
r10 18 65 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4480
+ $Y=0.1980 $X2=0.4300 $Y2=0.1980
r11 23 64 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1980 $X2=0.4590 $Y2=0.1765
r12 63 64 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1170 $X2=0.4590 $Y2=0.1765
r13 19 22 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0575 $X2=0.4590 $Y2=0.0360
r14 19 63 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0575 $X2=0.4590 $Y2=0.1170
r15 61 62 0.264706 $w=1.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3340 $Y=0.0725 $X2=0.3385 $Y2=0.0725
r16 3 61 0.705882 $w=1.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3220 $Y=0.0725 $X2=0.3340 $Y2=0.0725
r17 13 3 0.735294 $w=1.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0725 $X2=0.3220 $Y2=0.0725
r18 12 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0945 $X2=0.3220 $Y2=0.0945
r19 58 56 0.0675676 $w=3.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0455 $X2=0.3385 $Y2=0.0455
r20 3 56 0.391892 $w=3.7e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.0455 $X2=0.3385 $Y2=0.0455
r21 3 62 0.471383 $w=3.35517e-08 $l=3.06472e-08 $layer=N_src_drn
+ $thickness=1e-09 $X=0.3240 $Y=0.0455 $X2=0.3385 $Y2=0.0725
r22 11 3 0.391892 $w=3.7e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0455 $X2=0.3240 $Y2=0.0455
r23 57 11 0.0675676 $w=3.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0455 $X2=0.3095 $Y2=0.0455
r24 22 53 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4320 $Y2=0.0360
r25 3 46 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0540
+ $X2=0.3225 $Y2=0.0360
r26 52 53 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r27 51 52 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3800
+ $Y=0.0360 $X2=0.4050 $Y2=0.0360
r28 50 51 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3620
+ $Y=0.0360 $X2=0.3800 $Y2=0.0360
r29 49 50 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0360 $X2=0.3620 $Y2=0.0360
r30 48 49 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.0360 $X2=0.3510 $Y2=0.0360
r31 47 48 1.39914 $w=1.3e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.3315
+ $Y=0.0360 $X2=0.3375 $Y2=0.0360
r32 46 47 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3225
+ $Y=0.0360 $X2=0.3315 $Y2=0.0360
r33 45 46 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.3105
+ $Y=0.0360 $X2=0.3225 $Y2=0.0360
r34 44 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.3105 $Y2=0.0360
r35 43 44 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.2970 $Y2=0.0360
r36 42 43 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r37 41 42 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2180
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r38 40 41 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2000
+ $Y=0.0360 $X2=0.2180 $Y2=0.0360
r39 39 40 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.2000 $Y2=0.0360
r40 17 20 2.50689 $w=1.45385e-08 $l=1.86815e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1710 $Y=0.0360 $X2=0.1530 $Y2=0.0410
r41 17 39 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1710
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r42 20 37 3.32305 $w=1.42121e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1530 $Y=0.0410 $X2=0.1530 $Y2=0.0575
r43 36 37 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1530
+ $Y=0.0780 $X2=0.1530 $Y2=0.0575
r44 16 21 5.11339 $w=1.60414e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1530 $Y=0.1060 $X2=0.1530 $Y2=0.1350
r45 16 36 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1530
+ $Y=0.1060 $X2=0.1530 $Y2=0.0780
r46 21 34 3.01468 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1530
+ $Y=0.1350 $X2=0.1330 $Y2=0.1350
r47 10 30 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r48 33 34 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1195
+ $Y=0.1350 $X2=0.1330 $Y2=0.1350
r49 15 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1080 $Y=0.1350
+ $X2=0.1080 $Y2=0.1350
r50 15 33 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.1350 $X2=0.1195 $Y2=0.1350
r51 28 30 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1350 $X2=0.1350 $Y2=0.1350
r52 27 28 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1350 $X2=0.1225 $Y2=0.1350
r53 26 27 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1350 $X2=0.1080 $Y2=0.1350
r54 9 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r55 1 25 2.90696 $w=2.1681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0705 $Y2=0.1350
r56 1 26 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1350
r57 9 25 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.0810 $Y=0.1350 $X2=0.0705 $Y2=0.1350
r58 9 26 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1350
.ends


*
.SUBCKT AO32x2_ASAP7_75t_R VSS VDD A3 A2 A1 B1 B2 Y
*
* VSS VSS
* VDD VDD
* A3 A3
* A2 A2
* A1 A1
* B1 B1
* B2 B2
* Y Y
*
*

MM21 N_MM21_d N_MM21_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM21@2 N_MM21@2_d N_MM21@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM1_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM5_g N_MM0_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM13 N_MM13_d N_MM14_g N_MM13_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM18 N_MM18_d N_MM15_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM20 N_MM20_d N_MM21_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM20@2 N_MM20@2_d N_MM21@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1 N_MM1_d N_MM1_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM5_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM14 N_MM14_d N_MM14_g N_MM14_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM15 N_MM15_d N_MM15_g N_MM15_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2


*include "AO32x2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AO32x2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AO32x2_ASAP7_75t_R%NET26 VSS N_MM13_s N_MM18_d N_NET26_1
+ PM_AO32x2_ASAP7_75t_R%NET26
cc_1 N_NET26_1 N_MM14_g 0.0125199f
cc_2 N_NET26_1 N_MM15_g 0.0125836f
x_PM_AO32x2_ASAP7_75t_R%NET24 VSS N_MM2_d N_MM0_s N_NET24_1
+ PM_AO32x2_ASAP7_75t_R%NET24
cc_3 N_NET24_1 N_MM1_g 0.0173566f
cc_4 N_NET24_1 N_MM5_g 0.0173918f
x_PM_AO32x2_ASAP7_75t_R%NET25 VSS N_MM3_d N_MM2_s N_NET25_1
+ PM_AO32x2_ASAP7_75t_R%NET25
cc_5 N_NET25_1 N_MM3_g 0.0172674f
cc_6 N_NET25_1 N_MM1_g 0.017402f
x_PM_AO32x2_ASAP7_75t_R%A3 VSS A3 N_MM3_g N_A3_4 N_A3_1 PM_AO32x2_ASAP7_75t_R%A3
cc_7 N_A3_4 N_NET08_1 0.00093847f
cc_8 N_A3_4 N_NET08_17 0.00104187f
cc_9 N_A3_4 N_NET08_16 0.0024159f
cc_10 N_MM3_g N_MM21@2_g 0.00339575f
cc_11 N_A3_4 N_NET08_21 0.00718243f
x_PM_AO32x2_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_AO32x2_ASAP7_75t_R%noxref_16
cc_12 N_noxref_16_1 N_NET08_19 0.00094183f
cc_13 N_noxref_16_1 N_MM15_g 0.00369012f
x_PM_AO32x2_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_AO32x2_ASAP7_75t_R%noxref_17
cc_14 N_noxref_17_1 N_NET08_14 0.000919025f
cc_15 N_noxref_17_1 N_MM15_g 0.00366758f
cc_16 N_noxref_17_1 N_NET10_12 0.0266727f
cc_17 N_noxref_17_1 N_noxref_16_1 0.00205006f
x_PM_AO32x2_ASAP7_75t_R%A2 VSS A2 N_MM1_g N_A2_4 N_A2_1 PM_AO32x2_ASAP7_75t_R%A2
cc_18 N_A2_4 N_NET08_3 0.000273377f
cc_19 N_MM1_g N_NET08_12 0.000420151f
cc_20 N_A2_4 N_NET08_17 0.00147094f
cc_21 N_A2_4 N_NET08_21 0.00212953f
cc_22 N_A2_1 N_A3_1 0.00172449f
cc_23 N_A2_4 N_A3_4 0.00506546f
cc_24 N_MM1_g N_MM3_g 0.00838575f
x_PM_AO32x2_ASAP7_75t_R%B1 VSS B1 N_MM14_g N_B1_1 N_B1_4
+ PM_AO32x2_ASAP7_75t_R%B1
cc_25 N_MM14_g N_NET08_4 0.000725046f
cc_26 N_MM14_g N_NET08_12 0.00561202f
cc_27 N_MM14_g N_NET08_14 0.0112195f
cc_28 N_B1_1 N_NET08_3 0.000424207f
cc_29 N_B1_4 N_NET08_18 0.000585382f
cc_30 N_B1_1 N_NET08_11 0.00108447f
cc_31 N_B1_4 N_NET08_17 0.00128341f
cc_32 N_MM14_g N_NET08_3 0.00157594f
cc_33 N_B1_4 N_NET08_3 0.00247578f
cc_34 N_MM14_g N_NET08_11 0.0442257f
cc_35 N_B1_1 N_A1_1 0.00127224f
cc_36 N_B1_4 N_A1_4 0.00375689f
cc_37 N_MM14_g N_MM5_g 0.00668316f
x_PM_AO32x2_ASAP7_75t_R%B2 VSS B2 N_MM15_g N_B2_1 N_B2_4
+ PM_AO32x2_ASAP7_75t_R%B2
cc_38 N_MM15_g N_NET08_3 0.000256543f
cc_39 N_MM15_g N_NET08_4 0.00046712f
cc_40 N_B2_1 N_NET08_19 0.000619725f
cc_41 N_B2_1 N_NET08_14 0.000679797f
cc_42 N_B2_4 N_NET08_18 0.00115854f
cc_43 N_B2_4 N_NET08_17 0.00129383f
cc_44 N_B2_4 N_NET08_19 0.00637055f
cc_45 N_MM15_g N_NET08_14 0.0258981f
cc_46 N_B2_1 N_B1_1 0.00160927f
cc_47 N_B2_4 N_B1_4 0.00334114f
cc_48 N_MM15_g N_MM14_g 0.00968691f
x_PM_AO32x2_ASAP7_75t_R%A1 VSS A1 N_MM5_g N_A1_5 N_A1_1 N_A1_4
+ PM_AO32x2_ASAP7_75t_R%A1
cc_49 N_MM5_g N_NET08_11 0.0101542f
cc_50 N_MM5_g N_NET08_3 0.00188226f
cc_51 N_A1_5 N_NET08_18 0.000788256f
cc_52 N_A1_1 N_NET08_11 0.00081274f
cc_53 N_A1_4 N_NET08_17 0.00133392f
cc_54 N_A1_4 N_NET08_3 0.00200764f
cc_55 N_MM5_g N_NET08_12 0.0252683f
cc_56 N_MM5_g N_A2_1 0.00100157f
cc_57 N_A1_1 N_A2_1 0.00180131f
cc_58 N_A1_4 N_A2_4 0.00457536f
cc_59 N_MM5_g N_MM1_g 0.00760893f
x_PM_AO32x2_ASAP7_75t_R%NET10 VSS N_MM1_d N_MM4_d N_MM5_d N_MM14_s N_MM15_s
+ N_NET10_13 N_NET10_12 N_NET10_3 N_NET10_2 N_NET10_1 N_NET10_10 N_NET10_11
+ PM_AO32x2_ASAP7_75t_R%NET10
cc_60 N_NET10_13 N_NET08_14 0.00042508f
cc_61 N_NET10_13 N_NET08_19 0.000466248f
cc_62 N_NET10_12 N_NET08_14 0.00134789f
cc_63 N_NET10_3 N_NET08_18 0.000566851f
cc_64 N_NET10_13 N_NET08_23 0.000606249f
cc_65 N_NET10_13 N_NET08_4 0.000719911f
cc_66 N_NET10_2 N_NET08_4 0.000957994f
cc_67 N_NET10_3 N_NET08_4 0.0037906f
cc_68 N_NET10_13 N_NET08_18 0.00878776f
cc_69 N_NET10_1 N_MM3_g 0.000598865f
cc_70 N_NET10_1 N_A3_4 0.000964048f
cc_71 N_NET10_10 N_MM3_g 0.0252499f
cc_72 N_NET10_13 N_A2_4 0.00113015f
cc_73 N_NET10_1 N_A2_4 0.00143214f
cc_74 N_NET10_10 N_MM1_g 0.0256654f
cc_75 N_NET10_2 N_MM5_g 0.000863735f
cc_76 N_NET10_13 N_A1_5 0.00484616f
cc_77 N_NET10_11 N_MM5_g 0.025538f
cc_78 N_NET10_11 N_MM14_g 0.0255549f
cc_79 N_NET10_12 N_MM15_g 0.025616f
x_PM_AO32x2_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_AO32x2_ASAP7_75t_R%noxref_14
cc_80 N_noxref_14_1 N_MM21_g 0.00148339f
cc_81 N_noxref_14_1 N_Y_7 0.000755253f
x_PM_AO32x2_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_AO32x2_ASAP7_75t_R%noxref_15
cc_82 N_noxref_15_1 N_MM21_g 0.00147038f
cc_83 N_noxref_15_1 N_Y_8 0.000849689f
cc_84 N_noxref_15_1 N_noxref_14_1 0.00177626f
x_PM_AO32x2_ASAP7_75t_R%Y VSS Y N_MM21_d N_MM21@2_d N_MM20_d N_MM20@2_d N_Y_7
+ N_Y_9 N_Y_8 N_Y_14 N_Y_2 N_Y_1 PM_AO32x2_ASAP7_75t_R%Y
cc_85 N_Y_7 N_NET08_16 0.000354848f
cc_86 N_Y_7 N_NET08_15 0.000982539f
cc_87 N_Y_7 N_NET08_20 0.000451701f
cc_88 N_Y_7 N_NET08_1 0.0008826f
cc_89 N_Y_9 N_NET08_15 0.000908924f
cc_90 N_Y_8 N_MM21@2_g 0.0308509f
cc_91 N_Y_14 N_NET08_15 0.00157899f
cc_92 N_Y_2 N_MM21@2_g 0.00210948f
cc_93 N_Y_1 N_MM21@2_g 0.00211154f
cc_94 N_Y_14 N_NET08_16 0.00329032f
cc_95 N_Y_8 N_NET08_1 0.00452806f
cc_96 N_Y_7 N_MM21_g 0.0371568f
cc_97 N_Y_7 N_MM21@2_g 0.068582f
x_PM_AO32x2_ASAP7_75t_R%NET08 VSS N_MM21_g N_MM21@2_g N_MM0_d N_MM13_d N_MM14_d
+ N_MM15_d N_NET08_1 N_NET08_17 N_NET08_16 N_NET08_21 N_NET08_3 N_NET08_12
+ N_NET08_11 N_NET08_18 N_NET08_4 N_NET08_14 N_NET08_19 N_NET08_15 N_NET08_20
+ N_NET08_23 PM_AO32x2_ASAP7_75t_R%NET08
*END of AO32x2_ASAP7_75t_R.pxi
.ENDS
** Design:	AO331x1_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AO331x1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AO331x1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AO331x1_ASAP7_75t_R%NET32 VSS 2 3 1
c1 1 VSS 0.000990971f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3240 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3240 $Y2=0.0675
.ends

.subckt PM_AO331x1_ASAP7_75t_R%NET31 VSS 2 3 1
c1 1 VSS 0.000968743f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3780 $Y2=0.0675
.ends

.subckt PM_AO331x1_ASAP7_75t_R%N2 VSS 2 3 1
c1 1 VSS 0.00100671f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_AO331x1_ASAP7_75t_R%N1 VSS 2 3 1
c1 1 VSS 0.00101291f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2160 $Y2=0.0675
.ends

.subckt PM_AO331x1_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.00467662f
.ends

.subckt PM_AO331x1_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.00473277f
.ends

.subckt PM_AO331x1_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.00488656f
.ends

.subckt PM_AO331x1_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.00455837f
.ends

.subckt PM_AO331x1_ASAP7_75t_R%Y VSS 20 14 28 7 2 1 8 10 9
c1 1 VSS 0.00801092f
c2 2 VSS 0.00909286f
c3 7 VSS 0.00385734f
c4 8 VSS 0.0038338f
c5 9 VSS 0.00391753f
c6 10 VSS 0.00439325f
c7 11 VSS 0.00286075f
c8 12 VSS 0.00598222f
r1 28 27 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r2 8 27 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r3 2 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r4 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r5 12 23 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0270 $Y2=0.2125
r6 12 24 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0405 $Y2=0.2340
r7 22 23 8.51143 $w=1.3e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1760 $X2=0.0270 $Y2=0.2125
r8 21 22 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1500 $X2=0.0270 $Y2=0.1760
r9 20 21 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1475 $X2=0.0270 $Y2=0.1500
r10 20 19 9.91056 $w=1.3e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1475 $X2=0.0270 $Y2=0.1050
r11 9 11 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0540 $X2=0.0270 $Y2=0.0360
r12 9 19 11.8927 $w=1.3e-08 $l=5.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0540 $X2=0.0270 $Y2=0.1050
r13 10 15 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r14 10 11 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0405 $Y=0.0360 $X2=0.0270 $Y2=0.0360
r15 1 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0540 $Y2=0.0360
r16 14 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r17 7 13 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r18 2 8 1e-05
r19 1 7 1e-05
.ends

.subckt PM_AO331x1_ASAP7_75t_R%C VSS 6 3 1 4
c1 1 VSS 0.00809184f
c2 3 VSS 0.0453096f
c3 4 VSS 0.00482599f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1207 $X2=0.4590 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1150 $X2=0.4590 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1150 $X2=0.4590 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1350
+ $X2=0.4590 $Y2=0.1350
.ends

.subckt PM_AO331x1_ASAP7_75t_R%A2 VSS 8 3 4 1
c1 1 VSS 0.00635984f
c2 3 VSS 0.0463396f
c3 4 VSS 0.00466073f
r1 9 10 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1207 $X2=0.1890 $Y2=0.1350
r2 8 9 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1150 $X2=0.1890 $Y2=0.1207
r3 8 7 1.10765 $w=1.3e-08 $l=4.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1150 $X2=0.1890 $Y2=0.1102
r4 4 7 3.90593 $w=1.3e-08 $l=1.67e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0935 $X2=0.1890 $Y2=0.1102
r5 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r6 1 10 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AO331x1_ASAP7_75t_R%B2 VSS 6 3 4 1
c1 1 VSS 0.0072692f
c2 3 VSS 0.00984066f
c3 4 VSS 0.00475609f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1207 $X2=0.3510 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1150 $X2=0.3510 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1150 $X2=0.3510 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
.ends

.subckt PM_AO331x1_ASAP7_75t_R%A3 VSS 6 3 1 4
c1 1 VSS 0.00813583f
c2 3 VSS 0.0838473f
c3 4 VSS 0.00557256f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1207 $X2=0.1350 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1150 $X2=0.1350 $Y2=0.1207
r3 6 4 1.10765 $w=1.3e-08 $l=4.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1150 $X2=0.1350 $Y2=0.1102
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AO331x1_ASAP7_75t_R%A1 VSS 6 3 4 1
c1 1 VSS 0.00765577f
c2 3 VSS 0.0460661f
c3 4 VSS 0.00554335f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1207 $X2=0.2430 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1150 $X2=0.2430 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1150 $X2=0.2430 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AO331x1_ASAP7_75t_R%B1 VSS 6 3 1 4
c1 1 VSS 0.00776175f
c2 3 VSS 0.00914227f
c3 4 VSS 0.00495345f
r1 7 8 3.20636 $w=1.3e-08 $l=1.38e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1212 $X2=0.2970 $Y2=0.1350
r2 6 7 1.22425 $w=1.3e-08 $l=5.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1160 $X2=0.2970 $Y2=0.1212
r3 6 4 5.42166 $w=1.3e-08 $l=2.33e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1160 $X2=0.2970 $Y2=0.0927
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_AO331x1_ASAP7_75t_R%B3 VSS 6 3 4 1
c1 1 VSS 0.00870853f
c2 3 VSS 0.0470017f
c3 4 VSS 0.00516717f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1207 $X2=0.4050 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1150 $X2=0.4050 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1150 $X2=0.4050 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
.ends

.subckt PM_AO331x1_ASAP7_75t_R%NET24 VSS 12 13 25 26 2 8 9 1 7
c1 1 VSS 0.00292553f
c2 2 VSS 0.00318252f
c3 7 VSS 0.00214666f
c4 8 VSS 0.00219864f
c5 9 VSS 0.00236868f
r1 26 24 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r2 2 24 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r4 25 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r5 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.1980
r6 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4185
+ $Y=0.1980 $X2=0.4320 $Y2=0.1980
r7 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1980 $X2=0.4185 $Y2=0.1980
r8 18 19 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.3945
+ $Y=0.1980 $X2=0.4050 $Y2=0.1980
r9 17 18 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3765
+ $Y=0.1980 $X2=0.3945 $Y2=0.1980
r10 16 17 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1980 $X2=0.3765 $Y2=0.1980
r11 15 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.1980 $X2=0.3510 $Y2=0.1980
r12 14 15 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1980 $X2=0.3375 $Y2=0.1980
r13 9 14 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3115
+ $Y=0.1980 $X2=0.3240 $Y2=0.1980
r14 1 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.1980
r15 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r16 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r17 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r18 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
.ends

.subckt PM_AO331x1_ASAP7_75t_R%YB VSS 12 55 56 62 67 17 23 1 16 18 13 3 19 15 5
+ 4 20 14 21 24
c1 1 VSS 0.00372181f
c2 3 VSS 0.00590507f
c3 4 VSS 0.00814254f
c4 5 VSS 0.00560625f
c5 12 VSS 0.080121f
c6 13 VSS 0.00354944f
c7 14 VSS 0.00424343f
c8 15 VSS 0.00301828f
c9 16 VSS 0.00158536f
c10 17 VSS 0.00142542f
c11 18 VSS 0.000667489f
c12 19 VSS 0.0339995f
c13 20 VSS 0.00435393f
c14 21 VSS 0.000522543f
c15 22 VSS 0.00296417f
c16 23 VSS 0.000671647f
c17 24 VSS 0.00555042f
c18 25 VSS 0.00298279f
r1 15 5 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4840 $Y2=0.2025
r2 67 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r3 5 64 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2025
+ $X2=0.4860 $Y2=0.2340
r4 64 65 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.2340 $X2=0.4995 $Y2=0.2340
r5 24 60 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.2340 $X2=0.5130 $Y2=0.2160
r6 24 65 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.2340 $X2=0.4995 $Y2=0.2340
r7 14 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0675 $X2=0.4840 $Y2=0.0675
r8 62 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4715 $Y2=0.0675
r9 59 60 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1980 $X2=0.5130 $Y2=0.2160
r10 58 59 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1765 $X2=0.5130 $Y2=0.1980
r11 57 58 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1170 $X2=0.5130 $Y2=0.1765
r12 20 25 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.0575 $X2=0.5130 $Y2=0.0360
r13 20 57 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0575 $X2=0.5130 $Y2=0.1170
r14 56 54 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r15 3 54 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r16 13 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r17 55 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
r18 4 51 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0675
+ $X2=0.4860 $Y2=0.0360
r19 25 52 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.0360 $X2=0.4995 $Y2=0.0360
r20 3 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2700 $Y2=0.0360
r21 51 52 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.0360 $X2=0.4995 $Y2=0.0360
r22 50 51 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4740
+ $Y=0.0360 $X2=0.4860 $Y2=0.0360
r23 49 50 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4695
+ $Y=0.0360 $X2=0.4740 $Y2=0.0360
r24 48 49 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0360 $X2=0.4695 $Y2=0.0360
r25 47 48 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4485
+ $Y=0.0360 $X2=0.4590 $Y2=0.0360
r26 46 47 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4305
+ $Y=0.0360 $X2=0.4485 $Y2=0.0360
r27 45 46 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0360 $X2=0.4305 $Y2=0.0360
r28 44 45 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0360 $X2=0.4050 $Y2=0.0360
r29 43 44 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r30 42 43 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.3250
+ $Y=0.0360 $X2=0.3510 $Y2=0.0360
r31 41 42 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3070
+ $Y=0.0360 $X2=0.3250 $Y2=0.0360
r32 40 41 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.3070 $Y2=0.0360
r33 39 40 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2835
+ $Y=0.0360 $X2=0.2970 $Y2=0.0360
r34 38 39 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.2835 $Y2=0.0360
r35 37 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r36 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2565 $Y2=0.0360
r37 35 36 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r38 34 35 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r39 33 34 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.1630
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r40 19 22 0.682785 $w=1.75e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1450
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r41 19 33 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1450
+ $Y=0.0360 $X2=0.1630 $Y2=0.0360
r42 18 23 2.45586 $w=1.44e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.0540 $X2=0.1350 $Y2=0.0665
r43 18 22 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0540 $X2=0.1350 $Y2=0.0360
r44 17 21 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0720 $X2=0.0810 $Y2=0.0720
r45 17 23 4.55457 $w=1.3814e-08 $l=2.75545e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0720 $X2=0.1350 $Y2=0.0665
r46 21 31 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0720 $X2=0.0810 $Y2=0.0935
r47 16 29 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1160 $X2=0.0810 $Y2=0.1350
r48 16 31 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1160 $X2=0.0810 $Y2=0.0935
r49 12 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r50 1 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AO331x1_ASAP7_75t_R%NET034 VSS 16 17 33 34 37 38 1 10 13 2 11 12 3
c1 1 VSS 0.0100121f
c2 2 VSS 0.00700973f
c3 3 VSS 0.00447073f
c4 10 VSS 0.00452374f
c5 11 VSS 0.00332145f
c6 12 VSS 0.00212132f
c7 13 VSS 0.0223918f
r1 38 36 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r2 3 36 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r3 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3780 $Y2=0.2025
r4 37 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r5 34 32 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r6 2 32 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r7 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r8 33 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r9 3 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.2340
r10 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.2340
r11 28 29 9.211 $w=1.3e-08 $l=3.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.3385
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r12 27 28 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3070
+ $Y=0.2340 $X2=0.3385 $Y2=0.2340
r13 26 27 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.2340 $X2=0.3070 $Y2=0.2340
r14 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2835
+ $Y=0.2340 $X2=0.2970 $Y2=0.2340
r15 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.2835 $Y2=0.2340
r16 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r17 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2565 $Y2=0.2340
r18 21 22 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2430 $Y2=0.2340
r19 20 21 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r20 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1755
+ $Y=0.2340 $X2=0.1890 $Y2=0.2340
r21 18 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r22 13 18 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1495
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r23 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r24 16 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r25 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r26 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r27 17 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
.ends


*
.SUBCKT AO331x1_ASAP7_75t_R VSS VDD A3 A2 A1 B1 B2 B3 C Y
*
* VSS VSS
* VDD VDD
* A3 A3
* A2 A2
* A1 A1
* B1 B1
* B2 B2
* B3 B3
* C C
* Y Y
*
*

MM1 N_MM1_d N_MM1_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM16 N_MM16_d N_MM16_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM15 N_MM15_d N_MM25_g N_MM15_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM14 N_MM14_d N_MM24_g N_MM14_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM17 N_MM17_d N_MM20_g N_MM17_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM18 N_MM18_d N_MM21_g N_MM18_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM19 N_MM19_d N_MM23_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM22 N_MM22_d N_MM27_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM1_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM26 N_MM26_d N_MM16_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25 N_MM25_d N_MM25_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24 N_MM24_d N_MM24_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM20 N_MM20_d N_MM20_g N_MM20_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM21 N_MM21_d N_MM21_g N_MM21_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM23 N_MM23_d N_MM23_g N_MM23_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM27 N_MM27_d N_MM27_g N_MM27_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AO331x1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AO331x1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AO331x1_ASAP7_75t_R%NET32 VSS N_MM17_s N_MM18_d N_NET32_1
+ PM_AO331x1_ASAP7_75t_R%NET32
cc_1 N_NET32_1 N_MM20_g 0.0173032f
cc_2 N_NET32_1 N_MM21_g 0.0173936f
x_PM_AO331x1_ASAP7_75t_R%NET31 VSS N_MM18_s N_MM19_d N_NET31_1
+ PM_AO331x1_ASAP7_75t_R%NET31
cc_3 N_NET31_1 N_MM21_g 0.0173302f
cc_4 N_NET31_1 N_MM23_g 0.0173899f
x_PM_AO331x1_ASAP7_75t_R%N2 VSS N_MM16_d N_MM15_s N_N2_1
+ PM_AO331x1_ASAP7_75t_R%N2
cc_5 N_N2_1 N_MM16_g 0.0172756f
cc_6 N_N2_1 N_MM25_g 0.0174071f
x_PM_AO331x1_ASAP7_75t_R%N1 VSS N_MM15_d N_MM14_s N_N1_1
+ PM_AO331x1_ASAP7_75t_R%N1
cc_7 N_N1_1 N_MM25_g 0.0172906f
cc_8 N_N1_1 N_MM24_g 0.0173864f
x_PM_AO331x1_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_AO331x1_ASAP7_75t_R%noxref_19
cc_9 N_noxref_19_1 N_MM1_g 0.00146229f
cc_10 N_noxref_19_1 N_Y_8 0.0385647f
cc_11 N_noxref_19_1 N_noxref_18_1 0.00176553f
x_PM_AO331x1_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_AO331x1_ASAP7_75t_R%noxref_18
cc_12 N_noxref_18_1 N_MM1_g 0.00145369f
cc_13 N_noxref_18_1 N_Y_7 0.0384626f
x_PM_AO331x1_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_AO331x1_ASAP7_75t_R%noxref_20
cc_14 N_noxref_20_1 N_YB_20 0.000318238f
cc_15 N_noxref_20_1 N_YB_4 0.000505366f
cc_16 N_noxref_20_1 N_YB_14 0.0375276f
cc_17 N_noxref_20_1 N_MM27_g 0.0014503f
x_PM_AO331x1_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_AO331x1_ASAP7_75t_R%noxref_21
cc_18 N_noxref_21_1 N_YB_20 0.000318172f
cc_19 N_noxref_21_1 N_YB_5 0.000507441f
cc_20 N_noxref_21_1 N_YB_15 0.0377639f
cc_21 N_noxref_21_1 N_MM27_g 0.00144699f
cc_22 N_noxref_21_1 N_noxref_20_1 0.00176823f
x_PM_AO331x1_ASAP7_75t_R%Y VSS Y N_MM1_d N_MM0_d N_Y_7 N_Y_2 N_Y_1 N_Y_8 N_Y_10
+ N_Y_9 PM_AO331x1_ASAP7_75t_R%Y
cc_23 N_Y_7 N_YB_21 0.000223689f
cc_24 N_Y_7 N_YB_17 0.00039665f
cc_25 N_Y_7 N_YB_1 0.000785689f
cc_26 N_Y_2 N_MM1_g 0.00106757f
cc_27 N_Y_1 N_MM1_g 0.00143782f
cc_28 N_Y_8 N_YB_1 0.00165939f
cc_29 N_Y_10 N_YB_21 0.00265783f
cc_30 N_Y_9 N_YB_16 0.00459998f
cc_31 N_Y_8 N_MM1_g 0.015416f
cc_32 N_Y_7 N_MM1_g 0.0548551f
x_PM_AO331x1_ASAP7_75t_R%C VSS C N_MM27_g N_C_1 N_C_4 PM_AO331x1_ASAP7_75t_R%C
cc_33 N_MM27_g N_YB_15 0.0158971f
cc_34 N_C_1 N_YB_5 0.000815653f
cc_35 N_C_4 N_YB_19 0.00109537f
cc_36 N_MM27_g N_YB_5 0.00110236f
cc_37 N_MM27_g N_YB_4 0.00133751f
cc_38 N_C_1 N_YB_15 0.00171965f
cc_39 N_C_4 N_YB_20 0.00639089f
cc_40 N_MM27_g N_YB_14 0.0540039f
cc_41 N_MM27_g N_B3_1 0.000916468f
cc_42 N_C_4 N_B3_4 0.0032711f
cc_43 N_MM27_g N_MM23_g 0.00404287f
x_PM_AO331x1_ASAP7_75t_R%A2 VSS A2 N_MM25_g N_A2_4 N_A2_1
+ PM_AO331x1_ASAP7_75t_R%A2
cc_44 N_A2_4 N_YB_18 0.000136355f
cc_45 N_A2_4 N_YB_13 0.000145115f
cc_46 N_A2_4 N_YB_3 0.000268856f
cc_47 N_MM25_g N_YB_13 0.000457029f
cc_48 N_A2_4 N_YB_19 0.00133555f
cc_49 N_A2_4 N_YB_23 0.00280545f
cc_50 N_A2_1 N_A3_1 0.00133305f
cc_51 N_A2_4 N_A3_4 0.00379959f
cc_52 N_MM25_g N_MM16_g 0.00610095f
x_PM_AO331x1_ASAP7_75t_R%B2 VSS B2 N_MM21_g N_B2_4 N_B2_1
+ PM_AO331x1_ASAP7_75t_R%B2
cc_53 N_B2_4 N_YB_3 0.000269286f
cc_54 N_B2_4 N_YB_13 0.000415669f
cc_55 N_B2_4 N_YB_19 0.00332439f
cc_56 N_B2_1 N_B1_1 0.00126128f
cc_57 N_B2_4 N_B1_4 0.00343784f
cc_58 N_MM21_g N_MM20_g 0.00597422f
x_PM_AO331x1_ASAP7_75t_R%A3 VSS A3 N_MM16_g N_A3_1 N_A3_4
+ PM_AO331x1_ASAP7_75t_R%A3
cc_59 N_MM16_g N_YB_17 0.000362882f
cc_60 N_MM16_g N_YB_23 0.000548315f
cc_61 N_A3_1 N_YB_1 0.0019321f
cc_62 N_A3_4 N_YB_16 0.00337526f
cc_63 N_MM16_g N_MM1_g 0.00371803f
x_PM_AO331x1_ASAP7_75t_R%A1 VSS A1 N_MM24_g N_A1_4 N_A1_1
+ PM_AO331x1_ASAP7_75t_R%A1
cc_64 N_A1_4 N_YB_19 0.00129809f
cc_65 N_MM24_g N_YB_3 0.00154473f
cc_66 N_A1_4 N_YB_3 0.00197296f
cc_67 N_MM24_g N_YB_13 0.0365331f
cc_68 N_A1_1 N_A2_1 0.0012852f
cc_69 N_A1_4 N_A2_4 0.00460382f
cc_70 N_MM24_g N_MM25_g 0.00609516f
x_PM_AO331x1_ASAP7_75t_R%B1 VSS B1 N_MM20_g N_B1_1 N_B1_4
+ PM_AO331x1_ASAP7_75t_R%B1
cc_71 N_B1_1 N_YB_13 0.000842988f
cc_72 N_B1_4 N_YB_19 0.00130666f
cc_73 N_MM20_g N_YB_3 0.00154404f
cc_74 N_B1_4 N_YB_3 0.00176174f
cc_75 N_MM20_g N_YB_13 0.0357531f
cc_76 N_B1_1 N_A1_4 0.000836529f
cc_77 N_MM20_g N_MM24_g 0.0032795f
cc_78 N_B1_4 N_A1_4 0.00439129f
x_PM_AO331x1_ASAP7_75t_R%B3 VSS B3 N_MM23_g N_B3_4 N_B3_1
+ PM_AO331x1_ASAP7_75t_R%B3
cc_79 N_B3_4 N_YB_19 0.00335773f
cc_80 N_B3_1 N_B2_1 0.00141451f
cc_81 N_B3_4 N_B2_4 0.00358479f
cc_82 N_MM23_g N_MM21_g 0.00598122f
x_PM_AO331x1_ASAP7_75t_R%NET24 VSS N_MM20_d N_MM21_d N_MM23_d N_MM27_s
+ N_NET24_2 N_NET24_8 N_NET24_9 N_NET24_1 N_NET24_7 PM_AO331x1_ASAP7_75t_R%NET24
cc_83 N_NET24_2 N_YB_20 0.000372608f
cc_84 N_NET24_8 N_YB_15 0.0011152f
cc_85 N_NET24_9 N_YB_24 0.00133917f
cc_86 N_NET24_2 N_YB_5 0.00348718f
cc_87 N_NET24_9 N_B1_4 0.000612871f
cc_88 N_NET24_1 N_B1_4 0.000786663f
cc_89 N_NET24_1 N_MM20_g 0.00088404f
cc_90 N_NET24_7 N_MM20_g 0.033973f
cc_91 N_NET24_7 N_B2_1 0.000693955f
cc_92 N_NET24_1 N_MM21_g 0.000889588f
cc_93 N_NET24_9 N_B2_4 0.00120509f
cc_94 N_NET24_1 N_B2_4 0.00127174f
cc_95 N_NET24_7 N_MM21_g 0.0336264f
cc_96 N_NET24_2 N_MM23_g 0.000849808f
cc_97 N_NET24_8 N_B3_1 0.000860619f
cc_98 N_NET24_9 N_B3_4 0.00117636f
cc_99 N_NET24_2 N_B3_4 0.00131988f
cc_100 N_NET24_8 N_MM23_g 0.0336567f
cc_101 N_NET24_8 N_C_1 0.000686338f
cc_102 N_NET24_2 N_C_4 0.000763424f
cc_103 N_NET24_2 N_MM27_g 0.000865683f
cc_104 N_NET24_8 N_MM27_g 0.0341778f
cc_105 N_NET24_7 N_NET034_13 0.000554016f
cc_106 N_NET24_9 N_NET034_3 0.000681222f
cc_107 N_NET24_1 N_NET034_13 0.000771677f
cc_108 N_NET24_8 N_NET034_12 0.00111421f
cc_109 N_NET24_7 N_NET034_12 0.00111443f
cc_110 N_NET24_1 N_NET034_2 0.00133522f
cc_111 N_NET24_1 N_NET034_3 0.00274956f
cc_112 N_NET24_2 N_NET034_3 0.00424687f
cc_113 N_NET24_9 N_NET034_13 0.010197f
x_PM_AO331x1_ASAP7_75t_R%YB VSS N_MM1_g N_MM14_d N_MM17_d N_MM22_d N_MM27_d
+ N_YB_17 N_YB_23 N_YB_1 N_YB_16 N_YB_18 N_YB_13 N_YB_3 N_YB_19 N_YB_15 N_YB_5
+ N_YB_4 N_YB_20 N_YB_14 N_YB_21 N_YB_24 PM_AO331x1_ASAP7_75t_R%YB
x_PM_AO331x1_ASAP7_75t_R%NET034 VSS N_MM25_d N_MM26_d N_MM24_d N_MM20_s
+ N_MM21_s N_MM23_s N_NET034_1 N_NET034_10 N_NET034_13 N_NET034_2 N_NET034_11
+ N_NET034_12 N_NET034_3 PM_AO331x1_ASAP7_75t_R%NET034
cc_114 N_NET034_1 N_A3_4 0.00113226f
cc_115 N_NET034_1 N_MM16_g 0.00118095f
cc_116 N_NET034_10 N_MM16_g 0.0345543f
cc_117 N_NET034_10 N_A2_1 0.000650194f
cc_118 N_NET034_13 N_A2_4 0.00107078f
cc_119 N_NET034_1 N_MM25_g 0.00116257f
cc_120 N_NET034_1 N_A2_4 0.00161041f
cc_121 N_NET034_10 N_MM25_g 0.0334185f
cc_122 N_NET034_13 N_A1_4 0.00115944f
cc_123 N_NET034_2 N_MM24_g 0.00116329f
cc_124 N_NET034_2 N_A1_4 0.00165003f
cc_125 N_NET034_11 N_MM24_g 0.0340576f
cc_126 N_NET034_11 N_B1_1 0.00054468f
cc_127 N_NET034_2 N_MM20_g 0.000917773f
cc_128 N_NET034_11 N_MM20_g 0.033837f
cc_129 N_NET034_12 N_B2_1 0.000683578f
cc_130 N_NET034_3 N_MM21_g 0.000885284f
cc_131 N_NET034_12 N_MM21_g 0.0335386f
cc_132 N_NET034_12 N_B3_1 0.0007778f
cc_133 N_NET034_3 N_MM23_g 0.00087916f
cc_134 N_NET034_12 N_MM23_g 0.0334571f
*END of AO331x1_ASAP7_75t_R.pxi
.ENDS
** Design:	AO331x2_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AO331x2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AO331x2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AO331x2_ASAP7_75t_R%NET32 VSS 2 3 1
c1 1 VSS 0.000997736f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3780 $Y2=0.0675
.ends

.subckt PM_AO331x2_ASAP7_75t_R%NET31 VSS 2 3 1
c1 1 VSS 0.000963597f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4320 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4320 $Y2=0.0675
.ends

.subckt PM_AO331x2_ASAP7_75t_R%N2 VSS 2 3 1
c1 1 VSS 0.00101791f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2160 $Y2=0.0675
.ends

.subckt PM_AO331x2_ASAP7_75t_R%N1 VSS 2 3 1
c1 1 VSS 0.000994368f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2700 $Y2=0.0675
.ends

.subckt PM_AO331x2_ASAP7_75t_R%NET034 VSS 16 17 33 34 37 38 1 10 13 2 11 12 3
c1 1 VSS 0.0100485f
c2 2 VSS 0.00697118f
c3 3 VSS 0.00442898f
c4 10 VSS 0.00457749f
c5 11 VSS 0.00338198f
c6 12 VSS 0.0021738f
c7 13 VSS 0.0223938f
r1 38 36 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r2 3 36 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r3 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r4 37 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r5 34 32 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r6 2 32 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r7 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r8 33 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r9 3 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.2340
r10 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.2340
r11 28 29 9.211 $w=1.3e-08 $l=3.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.3925
+ $Y=0.2340 $X2=0.4320 $Y2=0.2340
r12 27 28 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3610
+ $Y=0.2340 $X2=0.3925 $Y2=0.2340
r13 26 27 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.2340 $X2=0.3610 $Y2=0.2340
r14 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.2340 $X2=0.3510 $Y2=0.2340
r15 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.2340 $X2=0.3375 $Y2=0.2340
r16 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3105
+ $Y=0.2340 $X2=0.3240 $Y2=0.2340
r17 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.2340 $X2=0.3105 $Y2=0.2340
r18 21 22 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.2970 $Y2=0.2340
r19 20 21 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r20 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.2340 $X2=0.2430 $Y2=0.2340
r21 18 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2295 $Y2=0.2340
r22 13 18 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2035
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r23 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.2340
r24 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r25 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r26 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r27 16 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
.ends

.subckt PM_AO331x2_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.0430745f
.ends

.subckt PM_AO331x2_ASAP7_75t_R%A1 VSS 6 3 1 4
c1 1 VSS 0.0076609f
c2 3 VSS 0.0460364f
c3 4 VSS 0.00550437f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1207 $X2=0.2970 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1150 $X2=0.2970 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1150 $X2=0.2970 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_AO331x2_ASAP7_75t_R%B2 VSS 6 3 4 1
c1 1 VSS 0.00744511f
c2 3 VSS 0.00986524f
c3 4 VSS 0.00483668f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1207 $X2=0.4050 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1150 $X2=0.4050 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1150 $X2=0.4050 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
.ends

.subckt PM_AO331x2_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.0430713f
.ends

.subckt PM_AO331x2_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.00475159f
.ends

.subckt PM_AO331x2_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.00467814f
.ends

.subckt PM_AO331x2_ASAP7_75t_R%Y VSS 22 15 16 31 32 7 8 9
c1 1 VSS 0.00977428f
c2 2 VSS 0.0109701f
c3 7 VSS 0.00468884f
c4 8 VSS 0.00467145f
c5 9 VSS 0.00770619f
c6 10 VSS 0.00438491f
c7 11 VSS 0.00343206f
c8 12 VSS 0.0063009f
r1 31 30 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r2 2 30 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r4 32 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
r5 2 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.2340
r6 26 27 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.2340 $X2=0.1080 $Y2=0.2340
r7 12 25 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.2340 $X2=0.0810 $Y2=0.2125
r8 12 26 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.2340 $X2=0.0945 $Y2=0.2340
r9 24 25 8.51143 $w=1.3e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1760 $X2=0.0810 $Y2=0.2125
r10 23 24 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1500 $X2=0.0810 $Y2=0.1760
r11 22 23 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1475 $X2=0.0810 $Y2=0.1500
r12 22 21 9.91056 $w=1.3e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1475 $X2=0.0810 $Y2=0.1050
r13 9 11 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0540 $X2=0.0810 $Y2=0.0360
r14 9 21 11.8927 $w=1.3e-08 $l=5.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0540 $X2=0.0810 $Y2=0.1050
r15 10 17 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.0360 $X2=0.1080 $Y2=0.0360
r16 10 11 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.0360 $X2=0.0810 $Y2=0.0360
r17 1 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1080 $Y2=0.0360
r18 16 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r19 1 14 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r20 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r21 15 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.0935 $Y2=0.0675
.ends

.subckt PM_AO331x2_ASAP7_75t_R%A3 VSS 6 3 1 4
c1 1 VSS 0.00786515f
c2 3 VSS 0.0835853f
c3 4 VSS 0.00539323f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1207 $X2=0.1890 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1150 $X2=0.1890 $Y2=0.1207
r3 6 4 1.10765 $w=1.3e-08 $l=4.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1150 $X2=0.1890 $Y2=0.1102
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AO331x2_ASAP7_75t_R%C VSS 6 3 1 4
c1 1 VSS 0.00795654f
c2 3 VSS 0.0453248f
c3 4 VSS 0.00486118f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1207 $X2=0.5130 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1150 $X2=0.5130 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1150 $X2=0.5130 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.1350
+ $X2=0.5130 $Y2=0.1350
.ends

.subckt PM_AO331x2_ASAP7_75t_R%A2 VSS 8 3 4 1
c1 1 VSS 0.00618775f
c2 3 VSS 0.0462924f
c3 4 VSS 0.00468052f
r1 9 10 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1207 $X2=0.2430 $Y2=0.1350
r2 8 9 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1150 $X2=0.2430 $Y2=0.1207
r3 8 7 1.10765 $w=1.3e-08 $l=4.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1150 $X2=0.2430 $Y2=0.1102
r4 4 7 3.90593 $w=1.3e-08 $l=1.67e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0935 $X2=0.2430 $Y2=0.1102
r5 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r6 1 10 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AO331x2_ASAP7_75t_R%B1 VSS 6 3 1 4
c1 1 VSS 0.00773996f
c2 3 VSS 0.00914948f
c3 4 VSS 0.00490145f
r1 7 8 3.20636 $w=1.3e-08 $l=1.38e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1212 $X2=0.3510 $Y2=0.1350
r2 6 7 1.22425 $w=1.3e-08 $l=5.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1160 $X2=0.3510 $Y2=0.1212
r3 6 4 5.42166 $w=1.3e-08 $l=2.33e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1160 $X2=0.3510 $Y2=0.0927
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
.ends

.subckt PM_AO331x2_ASAP7_75t_R%B3 VSS 6 3 4 1
c1 1 VSS 0.00827255f
c2 3 VSS 0.0467744f
c3 4 VSS 0.00494856f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1207 $X2=0.4590 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1150 $X2=0.4590 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1150 $X2=0.4590 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1350
+ $X2=0.4590 $Y2=0.1350
.ends

.subckt PM_AO331x2_ASAP7_75t_R%YB VSS 12 13 64 65 71 76 18 24 1 17 14 19 3 20
+ 15 16 5 4 21 23 22 25
c1 1 VSS 0.0077134f
c2 3 VSS 0.00602369f
c3 4 VSS 0.00849121f
c4 5 VSS 0.00594551f
c5 12 VSS 0.0807665f
c6 13 VSS 0.0805987f
c7 14 VSS 0.00525505f
c8 15 VSS 0.00605623f
c9 16 VSS 0.00484186f
c10 17 VSS 0.00217062f
c11 18 VSS 0.00159692f
c12 19 VSS 0.000671773f
c13 20 VSS 0.033654f
c14 21 VSS 0.00835638f
c15 22 VSS 0.000627341f
c16 23 VSS 0.00300404f
c17 24 VSS 0.000709787f
c18 25 VSS 0.00647611f
c19 26 VSS 0.00342605f
r1 16 5 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.2025 $X2=0.5380 $Y2=0.2025
r2 76 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.2025 $X2=0.5255 $Y2=0.2025
r3 5 73 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.2025
+ $X2=0.5400 $Y2=0.2340
r4 73 74 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.2340 $X2=0.5535 $Y2=0.2340
r5 25 69 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.2340 $X2=0.5670 $Y2=0.2160
r6 25 74 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.2340 $X2=0.5535 $Y2=0.2340
r7 15 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.0675 $X2=0.5380 $Y2=0.0675
r8 71 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.0675 $X2=0.5255 $Y2=0.0675
r9 68 69 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1980 $X2=0.5670 $Y2=0.2160
r10 67 68 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1765 $X2=0.5670 $Y2=0.1980
r11 66 67 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1170 $X2=0.5670 $Y2=0.1765
r12 21 26 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.0575 $X2=0.5670 $Y2=0.0360
r13 21 66 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0575 $X2=0.5670 $Y2=0.1170
r14 65 63 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r15 3 63 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r16 14 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3240 $Y2=0.0675
r17 64 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r18 4 60 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.0675
+ $X2=0.5400 $Y2=0.0360
r19 26 61 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.0360 $X2=0.5535 $Y2=0.0360
r20 3 47 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0675
+ $X2=0.3240 $Y2=0.0360
r21 60 61 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.0360 $X2=0.5535 $Y2=0.0360
r22 59 60 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.5280
+ $Y=0.0360 $X2=0.5400 $Y2=0.0360
r23 58 59 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.5235
+ $Y=0.0360 $X2=0.5280 $Y2=0.0360
r24 57 58 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0360 $X2=0.5235 $Y2=0.0360
r25 56 57 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.5025
+ $Y=0.0360 $X2=0.5130 $Y2=0.0360
r26 55 56 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4845
+ $Y=0.0360 $X2=0.5025 $Y2=0.0360
r27 54 55 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0360 $X2=0.4845 $Y2=0.0360
r28 53 54 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4590 $Y2=0.0360
r29 52 53 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r30 51 52 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.3790
+ $Y=0.0360 $X2=0.4050 $Y2=0.0360
r31 50 51 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3610
+ $Y=0.0360 $X2=0.3790 $Y2=0.0360
r32 49 50 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0360 $X2=0.3610 $Y2=0.0360
r33 48 49 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.0360 $X2=0.3510 $Y2=0.0360
r34 47 48 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.0360 $X2=0.3375 $Y2=0.0360
r35 46 47 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3105
+ $Y=0.0360 $X2=0.3240 $Y2=0.0360
r36 45 46 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.3105 $Y2=0.0360
r37 44 45 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.2970 $Y2=0.0360
r38 43 44 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r39 42 43 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2170
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r40 20 23 0.682785 $w=1.75e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1990
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r41 20 42 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1990
+ $Y=0.0360 $X2=0.2170 $Y2=0.0360
r42 19 24 2.45586 $w=1.44e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0540 $X2=0.1890 $Y2=0.0665
r43 19 23 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0540 $X2=0.1890 $Y2=0.0360
r44 18 22 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1620 $Y=0.0720 $X2=0.1350 $Y2=0.0720
r45 18 24 4.55457 $w=1.3814e-08 $l=2.75545e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1620 $Y=0.0720 $X2=0.1890 $Y2=0.0665
r46 22 40 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.0720 $X2=0.1350 $Y2=0.0935
r47 17 38 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1160 $X2=0.1350 $Y2=0.1350
r48 17 40 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1160 $X2=0.1350 $Y2=0.0935
r49 13 34 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1350 $Y2=0.1350
r50 34 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
r51 33 34 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1255
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r52 31 33 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1350 $X2=0.1255 $Y2=0.1350
r53 30 31 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1350 $X2=0.1225 $Y2=0.1350
r54 29 30 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1350 $X2=0.1080 $Y2=0.1350
r55 12 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r56 1 28 3.20232 $w=2.13909e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0700 $Y2=0.1350
r57 1 29 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1350
r58 12 28 0.905388 $w=2.07755e-07 $l=1.1e-08 $layer=LIG $thickness=5.52727e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0700 $Y2=0.1350
r59 12 29 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1350
.ends

.subckt PM_AO331x2_ASAP7_75t_R%NET24 VSS 12 13 25 26 2 8 9 1 7
c1 1 VSS 0.00289331f
c2 2 VSS 0.00318347f
c3 7 VSS 0.00212922f
c4 8 VSS 0.00217743f
c5 9 VSS 0.00218784f
r1 26 24 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r2 2 24 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4860 $Y2=0.2025
r4 25 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r5 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2025
+ $X2=0.4860 $Y2=0.1980
r6 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4725
+ $Y=0.1980 $X2=0.4860 $Y2=0.1980
r7 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1980 $X2=0.4725 $Y2=0.1980
r8 18 19 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4485
+ $Y=0.1980 $X2=0.4590 $Y2=0.1980
r9 17 18 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4305
+ $Y=0.1980 $X2=0.4485 $Y2=0.1980
r10 16 17 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1980 $X2=0.4305 $Y2=0.1980
r11 15 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3915
+ $Y=0.1980 $X2=0.4050 $Y2=0.1980
r12 14 15 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.1980 $X2=0.3915 $Y2=0.1980
r13 9 14 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3655
+ $Y=0.1980 $X2=0.3780 $Y2=0.1980
r14 1 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.1980
r15 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r16 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r17 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3780 $Y2=0.2025
r18 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
.ends


*
.SUBCKT AO331x2_ASAP7_75t_R VSS VDD A3 A2 A1 B1 B2 B3 C Y
*
* VSS VSS
* VDD VDD
* A3 A3
* A2 A2
* A1 A1
* B1 B1
* B2 B2
* B3 B3
* C C
* Y Y
*
*

MM1 N_MM1_d N_MM1_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1@2 N_MM1@2_d N_MM0@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM16 N_MM16_d N_MM26_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM15 N_MM15_d N_MM25_g N_MM15_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM14 N_MM14_d N_MM24_g N_MM14_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM17 N_MM17_d N_MM20_g N_MM17_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM18 N_MM18_d N_MM21_g N_MM18_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM19 N_MM19_d N_MM23_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM22 N_MM22_d N_MM27_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM1_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@2 N_MM0@2_d N_MM0@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM26 N_MM26_d N_MM26_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25 N_MM25_d N_MM25_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24 N_MM24_d N_MM24_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM20 N_MM20_d N_MM20_g N_MM20_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM21 N_MM21_d N_MM21_g N_MM21_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM23 N_MM23_d N_MM23_g N_MM23_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM27 N_MM27_d N_MM27_g N_MM27_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AO331x2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AO331x2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AO331x2_ASAP7_75t_R%NET32 VSS N_MM17_s N_MM18_d N_NET32_1
+ PM_AO331x2_ASAP7_75t_R%NET32
cc_1 N_NET32_1 N_MM20_g 0.0173794f
cc_2 N_NET32_1 N_MM21_g 0.0173111f
x_PM_AO331x2_ASAP7_75t_R%NET31 VSS N_MM18_s N_MM19_d N_NET31_1
+ PM_AO331x2_ASAP7_75t_R%NET31
cc_3 N_NET31_1 N_MM21_g 0.0174276f
cc_4 N_NET31_1 N_MM23_g 0.0172966f
x_PM_AO331x2_ASAP7_75t_R%N2 VSS N_MM16_d N_MM15_s N_N2_1
+ PM_AO331x2_ASAP7_75t_R%N2
cc_5 N_N2_1 N_MM26_g 0.0173529f
cc_6 N_N2_1 N_MM25_g 0.0173167f
x_PM_AO331x2_ASAP7_75t_R%N1 VSS N_MM15_d N_MM14_s N_N1_1
+ PM_AO331x2_ASAP7_75t_R%N1
cc_7 N_N1_1 N_MM25_g 0.0173922f
cc_8 N_N1_1 N_MM24_g 0.0173027f
x_PM_AO331x2_ASAP7_75t_R%NET034 VSS N_MM26_d N_MM25_d N_MM24_d N_MM20_s
+ N_MM21_s N_MM23_s N_NET034_1 N_NET034_10 N_NET034_13 N_NET034_2 N_NET034_11
+ N_NET034_12 N_NET034_3 PM_AO331x2_ASAP7_75t_R%NET034
cc_9 N_NET034_1 N_A3_4 0.00103248f
cc_10 N_NET034_1 N_MM26_g 0.0011798f
cc_11 N_NET034_10 N_MM26_g 0.0348497f
cc_12 N_NET034_10 N_A2_1 0.000668046f
cc_13 N_NET034_13 N_A2_4 0.00112343f
cc_14 N_NET034_1 N_MM25_g 0.00116916f
cc_15 N_NET034_1 N_A2_4 0.00155571f
cc_16 N_NET034_10 N_MM25_g 0.0335197f
cc_17 N_NET034_2 N_MM24_g 0.00118733f
cc_18 N_NET034_13 N_A1_4 0.00125221f
cc_19 N_NET034_2 N_A1_4 0.00164817f
cc_20 N_NET034_11 N_MM24_g 0.0343153f
cc_21 N_NET034_11 N_B1_1 0.000567289f
cc_22 N_NET034_2 N_MM20_g 0.000934164f
cc_23 N_NET034_11 N_MM20_g 0.0339604f
cc_24 N_NET034_12 N_B2_1 0.000646102f
cc_25 N_NET034_3 N_MM21_g 0.000892878f
cc_26 N_NET034_12 N_MM21_g 0.0338155f
cc_27 N_NET034_12 N_B3_1 0.000558959f
cc_28 N_NET034_3 N_MM23_g 0.00088391f
cc_29 N_NET034_12 N_MM23_g 0.0335526f
x_PM_AO331x2_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_AO331x2_ASAP7_75t_R%noxref_18
cc_30 N_noxref_18_1 N_MM1_g 0.00149989f
x_PM_AO331x2_ASAP7_75t_R%A1 VSS A1 N_MM24_g N_A1_1 N_A1_4
+ PM_AO331x2_ASAP7_75t_R%A1
cc_31 N_MM24_g N_YB_3 0.00182785f
cc_32 N_A1_1 N_YB_14 0.000890506f
cc_33 N_A1_4 N_YB_20 0.00128229f
cc_34 N_A1_4 N_YB_3 0.00195249f
cc_35 N_MM24_g N_YB_14 0.0356073f
cc_36 N_A1_1 N_A2_1 0.00134057f
cc_37 N_A1_4 N_A2_4 0.00458345f
cc_38 N_MM24_g N_MM25_g 0.00608886f
x_PM_AO331x2_ASAP7_75t_R%B2 VSS B2 N_MM21_g N_B2_4 N_B2_1
+ PM_AO331x2_ASAP7_75t_R%B2
cc_39 N_B2_4 N_YB_3 0.000268737f
cc_40 N_B2_4 N_YB_14 0.000417594f
cc_41 N_B2_4 N_YB_20 0.00324889f
cc_42 N_B2_1 N_B1_1 0.00132243f
cc_43 N_B2_4 N_B1_4 0.0034471f
cc_44 N_MM21_g N_MM20_g 0.00600733f
x_PM_AO331x2_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_AO331x2_ASAP7_75t_R%noxref_19
cc_45 N_noxref_19_1 N_MM1_g 0.00149397f
cc_46 N_noxref_19_1 N_noxref_18_1 0.00179775f
x_PM_AO331x2_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_AO331x2_ASAP7_75t_R%noxref_20
cc_47 N_noxref_20_1 N_YB_21 0.000326931f
cc_48 N_noxref_20_1 N_YB_4 0.000503912f
cc_49 N_noxref_20_1 N_YB_15 0.0376389f
cc_50 N_noxref_20_1 N_MM27_g 0.0014608f
x_PM_AO331x2_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_AO331x2_ASAP7_75t_R%noxref_21
cc_51 N_noxref_21_1 N_YB_21 0.000327027f
cc_52 N_noxref_21_1 N_YB_5 0.00050983f
cc_53 N_noxref_21_1 N_YB_16 0.0377463f
cc_54 N_noxref_21_1 N_MM27_g 0.00144766f
cc_55 N_noxref_21_1 N_noxref_20_1 0.00177257f
x_PM_AO331x2_ASAP7_75t_R%Y VSS Y N_MM1_d N_MM1@2_d N_MM0@2_d N_MM0_d N_Y_7
+ N_Y_8 N_Y_9 PM_AO331x2_ASAP7_75t_R%Y
cc_56 N_Y_7 N_YB_23 0.000153312f
cc_57 N_Y_7 N_YB_22 0.00280606f
cc_58 N_Y_7 N_YB_18 0.000395056f
cc_59 N_Y_7 N_YB_1 0.000644537f
cc_60 N_Y_8 N_YB_1 0.00490347f
cc_61 N_Y_9 N_YB_17 0.00502461f
cc_62 N_Y_8 N_MM1_g 0.0296319f
cc_63 N_Y_7 N_MM0@2_g 0.0365862f
cc_64 N_Y_7 N_MM1_g 0.0721255f
x_PM_AO331x2_ASAP7_75t_R%A3 VSS A3 N_MM26_g N_A3_1 N_A3_4
+ PM_AO331x2_ASAP7_75t_R%A3
cc_65 N_MM26_g N_YB_18 0.000357948f
cc_66 N_MM26_g N_YB_24 0.000628804f
cc_67 N_A3_1 N_YB_1 0.00188592f
cc_68 N_A3_4 N_YB_17 0.00319736f
cc_69 N_MM26_g N_MM0@2_g 0.00379353f
x_PM_AO331x2_ASAP7_75t_R%C VSS C N_MM27_g N_C_1 N_C_4 PM_AO331x2_ASAP7_75t_R%C
cc_70 N_MM27_g N_YB_16 0.0158853f
cc_71 N_C_1 N_YB_5 0.000840091f
cc_72 N_C_4 N_YB_20 0.00109617f
cc_73 N_MM27_g N_YB_5 0.00109978f
cc_74 N_MM27_g N_YB_4 0.00134091f
cc_75 N_C_1 N_YB_16 0.0016395f
cc_76 N_C_4 N_YB_21 0.00618706f
cc_77 N_MM27_g N_YB_15 0.0541194f
cc_78 N_MM27_g N_B3_1 0.000824848f
cc_79 N_C_4 N_B3_4 0.00314531f
cc_80 N_MM27_g N_MM23_g 0.00411447f
x_PM_AO331x2_ASAP7_75t_R%A2 VSS A2 N_MM25_g N_A2_4 N_A2_1
+ PM_AO331x2_ASAP7_75t_R%A2
cc_81 N_A2_4 N_YB_14 0.000252994f
cc_82 N_A2_4 N_YB_19 0.000136624f
cc_83 N_A2_4 N_YB_3 0.000268503f
cc_84 N_MM25_g N_YB_14 0.000470393f
cc_85 N_A2_4 N_YB_20 0.00131677f
cc_86 N_A2_4 N_YB_24 0.00276582f
cc_87 N_A2_1 N_A3_1 0.00135364f
cc_88 N_A2_4 N_A3_4 0.00377506f
cc_89 N_MM25_g N_MM26_g 0.00614298f
x_PM_AO331x2_ASAP7_75t_R%B1 VSS B1 N_MM20_g N_B1_1 N_B1_4
+ PM_AO331x2_ASAP7_75t_R%B1
cc_90 N_B1_1 N_YB_14 0.000889953f
cc_91 N_B1_4 N_YB_20 0.00129994f
cc_92 N_MM20_g N_YB_3 0.00156865f
cc_93 N_B1_4 N_YB_3 0.00181407f
cc_94 N_MM20_g N_YB_14 0.035654f
cc_95 N_B1_1 N_A1_4 0.00088641f
cc_96 N_MM20_g N_MM24_g 0.00327853f
cc_97 N_B1_4 N_A1_4 0.00447917f
x_PM_AO331x2_ASAP7_75t_R%B3 VSS B3 N_MM23_g N_B3_4 N_B3_1
+ PM_AO331x2_ASAP7_75t_R%B3
cc_98 N_B3_4 N_YB_15 0.00016895f
cc_99 N_B3_4 N_YB_20 0.00312375f
cc_100 N_B3_1 N_B2_1 0.00131701f
cc_101 N_B3_4 N_B2_4 0.00338503f
cc_102 N_MM23_g N_MM21_g 0.00597838f
x_PM_AO331x2_ASAP7_75t_R%YB VSS N_MM1_g N_MM0@2_g N_MM14_d N_MM17_d N_MM22_d
+ N_MM27_d N_YB_18 N_YB_24 N_YB_1 N_YB_17 N_YB_14 N_YB_19 N_YB_3 N_YB_20
+ N_YB_15 N_YB_16 N_YB_5 N_YB_4 N_YB_21 N_YB_23 N_YB_22 N_YB_25
+ PM_AO331x2_ASAP7_75t_R%YB
x_PM_AO331x2_ASAP7_75t_R%NET24 VSS N_MM20_d N_MM21_d N_MM23_d N_MM27_s
+ N_NET24_2 N_NET24_8 N_NET24_9 N_NET24_1 N_NET24_7 PM_AO331x2_ASAP7_75t_R%NET24
cc_103 N_NET24_2 N_YB_21 0.000387955f
cc_104 N_NET24_8 N_YB_16 0.0011068f
cc_105 N_NET24_9 N_YB_25 0.00124604f
cc_106 N_NET24_2 N_YB_5 0.00347834f
cc_107 N_NET24_9 N_B1_4 0.000602231f
cc_108 N_NET24_1 N_B1_4 0.000731744f
cc_109 N_NET24_1 N_MM20_g 0.000885352f
cc_110 N_NET24_7 N_MM20_g 0.0338746f
cc_111 N_NET24_7 N_B2_1 0.000730937f
cc_112 N_NET24_1 N_MM21_g 0.000877593f
cc_113 N_NET24_9 N_B2_4 0.00110756f
cc_114 N_NET24_1 N_B2_4 0.00121385f
cc_115 N_NET24_7 N_MM21_g 0.0333829f
cc_116 N_NET24_8 N_B3_1 0.000591108f
cc_117 N_NET24_2 N_MM23_g 0.000843672f
cc_118 N_NET24_9 N_B3_4 0.00110701f
cc_119 N_NET24_2 N_B3_4 0.00121631f
cc_120 N_NET24_8 N_MM23_g 0.0335105f
cc_121 N_NET24_8 N_C_1 0.000692853f
cc_122 N_NET24_2 N_C_4 0.000739528f
cc_123 N_NET24_2 N_MM27_g 0.000862829f
cc_124 N_NET24_8 N_MM27_g 0.033976f
cc_125 N_NET24_7 N_NET034_13 0.000552738f
cc_126 N_NET24_9 N_NET034_3 0.000666108f
cc_127 N_NET24_1 N_NET034_13 0.000698446f
cc_128 N_NET24_7 N_NET034_11 0.00111162f
cc_129 N_NET24_7 N_NET034_12 0.00111192f
cc_130 N_NET24_2 N_NET034_3 0.00121563f
cc_131 N_NET24_1 N_NET034_3 0.00302384f
cc_132 N_NET24_1 N_NET034_2 0.00407046f
cc_133 N_NET24_9 N_NET034_13 0.00977738f
*END of AO331x2_ASAP7_75t_R.pxi
.ENDS
** Design:	AO332x1_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AO332x1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AO332x1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AO332x1_ASAP7_75t_R%NET061 VSS 2 3 1
c1 1 VSS 0.00102077f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4860 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0675 $X2=0.4860 $Y2=0.0675
.ends

.subckt PM_AO332x1_ASAP7_75t_R%NET063 VSS 2 3 1
c1 1 VSS 0.000970755f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3240 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3240 $Y2=0.0675
.ends

.subckt PM_AO332x1_ASAP7_75t_R%NET25 VSS 2 3 1
c1 1 VSS 0.000973405f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_AO332x1_ASAP7_75t_R%NET064 VSS 2 3 1
c1 1 VSS 0.000984958f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3780 $Y2=0.0675
.ends

.subckt PM_AO332x1_ASAP7_75t_R%NET26 VSS 2 3 1
c1 1 VSS 0.000962031f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2160 $Y2=0.0675
.ends

.subckt PM_AO332x1_ASAP7_75t_R%NET031 VSS 20 21 38 39 42 43 10 1 13 11 2 15 12 3
c1 1 VSS 0.0100716f
c2 2 VSS 0.00558338f
c3 3 VSS 0.00309579f
c4 10 VSS 0.00451746f
c5 11 VSS 0.00333873f
c6 12 VSS 0.00213955f
c7 13 VSS 0.00836819f
c8 14 VSS 0.000550778f
c9 15 VSS 0.00183748f
c10 16 VSS 0.000577327f
c11 17 VSS 0.00264588f
r1 43 41 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r2 3 41 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r3 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3780 $Y2=0.2025
r4 42 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r5 39 37 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r6 2 37 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r7 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r8 38 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r9 3 34 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.1980
r10 2 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.1980
r11 33 34 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3645
+ $Y=0.1980 $X2=0.3780 $Y2=0.1980
r12 32 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1980 $X2=0.3645 $Y2=0.1980
r13 31 32 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.3250
+ $Y=0.1980 $X2=0.3510 $Y2=0.1980
r14 30 31 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3070
+ $Y=0.1980 $X2=0.3250 $Y2=0.1980
r15 29 30 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1980 $X2=0.3070 $Y2=0.1980
r16 28 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2835
+ $Y=0.1980 $X2=0.2970 $Y2=0.1980
r17 27 28 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1980 $X2=0.2835 $Y2=0.1980
r18 15 27 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.1980 $X2=0.2700 $Y2=0.1980
r19 15 16 1.40651 $w=1.51875e-08 $l=1.45774e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2565 $Y=0.1980 $X2=0.2430 $Y2=0.2035
r20 14 17 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2160 $X2=0.2430 $Y2=0.2340
r21 14 16 2.45586 $w=1.44e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.2160 $X2=0.2430 $Y2=0.2035
r22 17 25 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.2340 $X2=0.2160 $Y2=0.2340
r23 24 25 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r24 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1755
+ $Y=0.2340 $X2=0.1890 $Y2=0.2340
r25 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r26 13 22 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1495
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r27 1 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r28 21 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r29 1 19 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r30 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r31 20 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
.ends

.subckt PM_AO332x1_ASAP7_75t_R%A3 VSS 6 3 1 4
c1 1 VSS 0.0078774f
c2 3 VSS 0.0837381f
c3 4 VSS 0.0055009f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1207 $X2=0.1350 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1150 $X2=0.1350 $Y2=0.1207
r3 6 4 1.10765 $w=1.3e-08 $l=4.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1150 $X2=0.1350 $Y2=0.1102
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AO332x1_ASAP7_75t_R%A2 VSS 6 3 4 1
c1 1 VSS 0.00646905f
c2 3 VSS 0.0464264f
c3 4 VSS 0.00490296f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1207 $X2=0.1890 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1150 $X2=0.1890 $Y2=0.1207
r3 6 4 1.10765 $w=1.3e-08 $l=4.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1150 $X2=0.1890 $Y2=0.1102
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AO332x1_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.00466082f
.ends

.subckt PM_AO332x1_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.0047668f
.ends

.subckt PM_AO332x1_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.00475751f
.ends

.subckt PM_AO332x1_ASAP7_75t_R%C2 VSS 6 3 4 1
c1 1 VSS 0.00691936f
c2 3 VSS 0.0463514f
c3 4 VSS 0.00470529f
r1 7 8 3.43955 $w=1.3e-08 $l=1.48e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1202 $X2=0.4590 $Y2=0.1350
r2 6 7 1.45744 $w=1.3e-08 $l=6.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1140 $X2=0.4590 $Y2=0.1202
r3 6 4 5.18847 $w=1.3e-08 $l=2.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1140 $X2=0.4590 $Y2=0.0917
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1350
+ $X2=0.4590 $Y2=0.1350
.ends

.subckt PM_AO332x1_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.00608609f
.ends

.subckt PM_AO332x1_ASAP7_75t_R%B1 VSS 6 3 1 4
c1 1 VSS 0.0077788f
c2 3 VSS 0.00916332f
c3 4 VSS 0.0049004f
r1 7 8 3.20636 $w=1.3e-08 $l=1.38e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1212 $X2=0.2970 $Y2=0.1350
r2 6 7 1.22425 $w=1.3e-08 $l=5.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1160 $X2=0.2970 $Y2=0.1212
r3 6 4 5.42166 $w=1.3e-08 $l=2.33e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1160 $X2=0.2970 $Y2=0.0927
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_AO332x1_ASAP7_75t_R%B3 VSS 6 3 4 1
c1 1 VSS 0.00808861f
c2 3 VSS 0.0468375f
c3 4 VSS 0.00508659f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1207 $X2=0.4050 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1150 $X2=0.4050 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1150 $X2=0.4050 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
.ends

.subckt PM_AO332x1_ASAP7_75t_R%Y VSS 20 14 28 7 2 1 8 10 9
c1 1 VSS 0.00798591f
c2 2 VSS 0.00877959f
c3 7 VSS 0.00383944f
c4 8 VSS 0.00382936f
c5 9 VSS 0.00408422f
c6 10 VSS 0.00607498f
c7 11 VSS 0.00281047f
c8 12 VSS 0.0076565f
r1 28 27 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r2 8 27 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r3 2 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r4 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r5 12 23 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0270 $Y2=0.2125
r6 12 24 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0405 $Y2=0.2340
r7 22 23 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1755 $X2=0.0270 $Y2=0.2125
r8 21 22 6.99569 $w=1.3e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1455 $X2=0.0270 $Y2=0.1755
r9 20 21 1.39914 $w=1.3e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1395 $X2=0.0270 $Y2=0.1455
r10 20 19 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1395 $X2=0.0270 $Y2=0.1010
r11 9 11 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0540 $X2=0.0270 $Y2=0.0360
r12 9 19 10.9599 $w=1.3e-08 $l=4.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0540 $X2=0.0270 $Y2=0.1010
r13 10 15 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r14 10 11 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0405 $Y=0.0360 $X2=0.0270 $Y2=0.0360
r15 1 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0540 $Y2=0.0360
r16 14 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r17 7 13 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r18 2 8 1e-05
r19 1 7 1e-05
.ends

.subckt PM_AO332x1_ASAP7_75t_R%C1 VSS 6 3 1 4
c1 1 VSS 0.00692823f
c2 3 VSS 0.00864116f
c3 4 VSS 0.00433882f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1207 $X2=0.5130 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1150 $X2=0.5130 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1150 $X2=0.5130 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.1350
+ $X2=0.5130 $Y2=0.1350
.ends

.subckt PM_AO332x1_ASAP7_75t_R%A1 VSS 6 3 1 4
c1 1 VSS 0.00720477f
c2 3 VSS 0.0458769f
c3 4 VSS 0.00402147f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1207 $X2=0.2430 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1150 $X2=0.2430 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1150 $X2=0.2430 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AO332x1_ASAP7_75t_R%B2 VSS 6 3 4 1
c1 1 VSS 0.00741386f
c2 3 VSS 0.00987809f
c3 4 VSS 0.00487177f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1207 $X2=0.3510 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1150 $X2=0.3510 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1150 $X2=0.3510 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
.ends

.subckt PM_AO332x1_ASAP7_75t_R%NET018 VSS 12 56 57 61 69 70 17 24 1 16 13 18 3
+ 19 5 4 20 15 14 21 22 23 26
c1 1 VSS 0.00354107f
c2 3 VSS 0.00577217f
c3 4 VSS 0.00300248f
c4 5 VSS 0.00583248f
c5 12 VSS 0.080021f
c6 13 VSS 0.00322483f
c7 14 VSS 0.00306764f
c8 15 VSS 0.00251317f
c9 16 VSS 0.00148445f
c10 17 VSS 0.00128547f
c11 18 VSS 0.000654402f
c12 19 VSS 0.0382705f
c13 20 VSS 0.000841668f
c14 21 VSS 0.00260666f
c15 22 VSS 0.000458078f
c16 23 VSS 0.00285804f
c17 24 VSS 0.000638966f
c18 25 VSS 0.00285347f
c19 26 VSS 0.000886268f
r1 70 68 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r2 4 68 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r3 15 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4860 $Y2=0.2025
r4 69 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r5 4 65 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2025
+ $X2=0.4860 $Y2=0.1980
r6 65 66 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.1980 $X2=0.4995 $Y2=0.1980
r7 63 66 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1980 $X2=0.4995 $Y2=0.1980
r8 62 63 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.5390
+ $Y=0.1980 $X2=0.5130 $Y2=0.1980
r9 20 26 0.682785 $w=1.75e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5570
+ $Y=0.1980 $X2=0.5670 $Y2=0.1980
r10 20 62 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5570
+ $Y=0.1980 $X2=0.5390 $Y2=0.1980
r11 26 59 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.1980 $X2=0.5670 $Y2=0.1765
r12 14 5 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.0675 $X2=0.5380 $Y2=0.0675
r13 61 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.0675 $X2=0.5255 $Y2=0.0675
r14 58 59 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1170 $X2=0.5670 $Y2=0.1765
r15 21 25 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.0575 $X2=0.5670 $Y2=0.0360
r16 21 58 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0575 $X2=0.5670 $Y2=0.1170
r17 57 55 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r18 3 55 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r19 13 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r20 56 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
r21 5 52 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.0675
+ $X2=0.5400 $Y2=0.0360
r22 25 53 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.0360 $X2=0.5535 $Y2=0.0360
r23 3 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2700 $Y2=0.0360
r24 52 53 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.0360 $X2=0.5535 $Y2=0.0360
r25 51 52 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5265
+ $Y=0.0360 $X2=0.5400 $Y2=0.0360
r26 50 51 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0360 $X2=0.5265 $Y2=0.0360
r27 49 50 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.4875
+ $Y=0.0360 $X2=0.5130 $Y2=0.0360
r28 48 49 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4695
+ $Y=0.0360 $X2=0.4875 $Y2=0.0360
r29 47 48 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0360 $X2=0.4695 $Y2=0.0360
r30 46 47 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4590 $Y2=0.0360
r31 45 46 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r32 44 45 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.3945
+ $Y=0.0360 $X2=0.4050 $Y2=0.0360
r33 43 44 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3765
+ $Y=0.0360 $X2=0.3945 $Y2=0.0360
r34 42 43 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0360 $X2=0.3765 $Y2=0.0360
r35 41 42 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.0360 $X2=0.3510 $Y2=0.0360
r36 40 41 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.3240 $Y2=0.0360
r37 39 40 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2835
+ $Y=0.0360 $X2=0.2970 $Y2=0.0360
r38 38 39 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.2835 $Y2=0.0360
r39 37 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r40 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2565 $Y2=0.0360
r41 35 36 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r42 34 35 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r43 33 34 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.1630
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r44 19 23 0.682785 $w=1.75e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1450
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r45 19 33 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1450
+ $Y=0.0360 $X2=0.1630 $Y2=0.0360
r46 18 24 2.45586 $w=1.44e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.0540 $X2=0.1350 $Y2=0.0665
r47 18 23 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0540 $X2=0.1350 $Y2=0.0360
r48 24 31 4.08819 $w=1.38974e-08 $l=2.55979e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.0665 $X2=0.1100 $Y2=0.0720
r49 17 22 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0920 $Y=0.0720 $X2=0.0810 $Y2=0.0720
r50 17 31 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0920
+ $Y=0.0720 $X2=0.1100 $Y2=0.0720
r51 22 30 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0720 $X2=0.0810 $Y2=0.0935
r52 16 28 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1160 $X2=0.0810 $Y2=0.1350
r53 16 30 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1160 $X2=0.0810 $Y2=0.0935
r54 12 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r55 1 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AO332x1_ASAP7_75t_R%NET030 VSS 16 17 32 33 35 13 3 12 2 10 1 11
c1 1 VSS 0.00466381f
c2 2 VSS 0.00461712f
c3 3 VSS 0.00518943f
c4 10 VSS 0.00220499f
c5 11 VSS 0.00219791f
c6 12 VSS 0.0022606f
c7 13 VSS 0.0227354f
r1 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.2025 $X2=0.5380 $Y2=0.2025
r2 35 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.2025 $X2=0.5255 $Y2=0.2025
r3 33 31 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r4 2 31 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r5 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r6 32 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r7 3 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.2025
+ $X2=0.5400 $Y2=0.2340
r8 2 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.2340
r9 27 28 9.0944 $w=1.3e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.5010
+ $Y=0.2340 $X2=0.5400 $Y2=0.2340
r10 26 27 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4695
+ $Y=0.2340 $X2=0.5010 $Y2=0.2340
r11 25 26 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4695 $Y2=0.2340
r12 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4455
+ $Y=0.2340 $X2=0.4590 $Y2=0.2340
r13 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4455 $Y2=0.2340
r14 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4185
+ $Y=0.2340 $X2=0.4320 $Y2=0.2340
r15 21 22 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.2340 $X2=0.4185 $Y2=0.2340
r16 20 21 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.3945
+ $Y=0.2340 $X2=0.4050 $Y2=0.2340
r17 19 20 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3630
+ $Y=0.2340 $X2=0.3945 $Y2=0.2340
r18 18 19 9.0944 $w=1.3e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.2340 $X2=0.3630 $Y2=0.2340
r19 13 18 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3115
+ $Y=0.2340 $X2=0.3240 $Y2=0.2340
r20 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.2340
r21 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r22 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r23 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r24 16 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
.ends


*
.SUBCKT AO332x1_ASAP7_75t_R VSS VDD A3 A2 A1 B1 B2 B3 C2 C1 Y
*
* VSS VSS
* VDD VDD
* A3 A3
* A2 A2
* A1 A1
* B1 B1
* B2 B2
* B3 B3
* C2 C2
* C1 C1
* Y Y
*
*

MM13 N_MM13_d N_MM13_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM8_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM14 N_MM14_d N_MM9_g N_MM14_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM12 N_MM12_d N_MM6_g N_MM12_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 N_MM11_d N_MM5_g N_MM11_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM16 N_MM16_d N_MM0_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM17 N_MM17_d N_MM1_g N_MM17_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM15 N_MM15_d N_MM13_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM8_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM6_g N_MM6_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g N_MM4_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM0_g N_MM0_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AO332x1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AO332x1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AO332x1_ASAP7_75t_R%NET061 VSS N_MM16_d N_MM17_s N_NET061_1
+ PM_AO332x1_ASAP7_75t_R%NET061
cc_1 N_NET061_1 N_MM0_g 0.017335f
cc_2 N_NET061_1 N_MM1_g 0.0174454f
x_PM_AO332x1_ASAP7_75t_R%NET063 VSS N_MM12_s N_MM11_d N_NET063_1
+ PM_AO332x1_ASAP7_75t_R%NET063
cc_3 N_NET063_1 N_MM6_g 0.017225f
cc_4 N_NET063_1 N_MM5_g 0.0173651f
x_PM_AO332x1_ASAP7_75t_R%NET25 VSS N_MM3_d N_MM2_s N_NET25_1
+ PM_AO332x1_ASAP7_75t_R%NET25
cc_5 N_NET25_1 N_MM7_g 0.0172763f
cc_6 N_NET25_1 N_MM8_g 0.0174241f
x_PM_AO332x1_ASAP7_75t_R%NET064 VSS N_MM11_s N_MM10_d N_NET064_1
+ PM_AO332x1_ASAP7_75t_R%NET064
cc_7 N_NET064_1 N_MM5_g 0.0173406f
cc_8 N_NET064_1 N_MM4_g 0.0173473f
x_PM_AO332x1_ASAP7_75t_R%NET26 VSS N_MM2_d N_MM14_s N_NET26_1
+ PM_AO332x1_ASAP7_75t_R%NET26
cc_9 N_NET26_1 N_MM8_g 0.0172619f
cc_10 N_NET26_1 N_MM9_g 0.0173383f
x_PM_AO332x1_ASAP7_75t_R%NET031 VSS N_MM7_d N_MM8_d N_MM9_d N_MM6_s N_MM5_s
+ N_MM4_s N_NET031_10 N_NET031_1 N_NET031_13 N_NET031_11 N_NET031_2 N_NET031_15
+ N_NET031_12 N_NET031_3 PM_AO332x1_ASAP7_75t_R%NET031
cc_11 N_NET031_10 N_A3_1 0.00077317f
cc_12 N_NET031_1 N_A3_4 0.00111594f
cc_13 N_NET031_1 N_MM7_g 0.0011587f
cc_14 N_NET031_10 N_MM7_g 0.0339579f
cc_15 N_NET031_10 N_A2_1 0.000647654f
cc_16 N_NET031_13 N_A2_4 0.00100875f
cc_17 N_NET031_1 N_MM8_g 0.00114378f
cc_18 N_NET031_1 N_A2_4 0.00196951f
cc_19 N_NET031_10 N_MM8_g 0.0342042f
cc_20 N_NET031_11 N_A1_4 0.000470017f
cc_21 N_NET031_11 N_A1_1 0.000672334f
cc_22 N_NET031_2 N_MM9_g 0.000881893f
cc_23 N_NET031_2 N_A1_4 0.00108461f
cc_24 N_NET031_11 N_MM9_g 0.0340457f
cc_25 N_NET031_11 N_B1_1 0.000616959f
cc_26 N_NET031_2 N_MM6_g 0.000876696f
cc_27 N_NET031_15 N_B1_4 0.00113657f
cc_28 N_NET031_2 N_B1_4 0.00125444f
cc_29 N_NET031_11 N_MM6_g 0.0336777f
cc_30 N_NET031_12 N_B2_1 0.000817576f
cc_31 N_NET031_3 N_MM5_g 0.00086063f
cc_32 N_NET031_15 N_B2_4 0.00114262f
cc_33 N_NET031_3 N_B2_4 0.00122286f
cc_34 N_NET031_12 N_MM5_g 0.033643f
cc_35 N_NET031_12 N_B3_4 0.000573728f
cc_36 N_NET031_12 N_B3_1 0.000739774f
cc_37 N_NET031_3 N_B3_4 0.000758694f
cc_38 N_NET031_3 N_MM4_g 0.000865311f
cc_39 N_NET031_12 N_MM4_g 0.0335356f
x_PM_AO332x1_ASAP7_75t_R%A3 VSS A3 N_MM7_g N_A3_1 N_A3_4
+ PM_AO332x1_ASAP7_75t_R%A3
cc_40 N_MM7_g N_NET018_17 0.000444474f
cc_41 N_MM7_g N_NET018_24 0.000469781f
cc_42 N_MM7_g N_NET018_1 0.000846414f
cc_43 N_A3_1 N_NET018_1 0.000970247f
cc_44 N_A3_4 N_NET018_16 0.00319942f
cc_45 N_MM7_g N_MM13_g 0.00375405f
x_PM_AO332x1_ASAP7_75t_R%A2 VSS A2 N_MM8_g N_A2_4 N_A2_1
+ PM_AO332x1_ASAP7_75t_R%A2
cc_46 N_A2_4 N_NET018_13 0.00024788f
cc_47 N_A2_4 N_NET018_18 0.000188886f
cc_48 N_A2_4 N_NET018_3 0.000278616f
cc_49 N_MM8_g N_NET018_13 0.000454535f
cc_50 N_A2_4 N_NET018_19 0.00130209f
cc_51 N_A2_4 N_NET018_24 0.00285763f
cc_52 N_A2_1 N_A3_1 0.00131305f
cc_53 N_A2_4 N_A3_4 0.00392067f
cc_54 N_MM8_g N_MM7_g 0.00605292f
x_PM_AO332x1_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_AO332x1_ASAP7_75t_R%noxref_20
cc_55 N_noxref_20_1 N_MM13_g 0.00145516f
cc_56 N_noxref_20_1 N_Y_7 0.0385931f
x_PM_AO332x1_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_AO332x1_ASAP7_75t_R%noxref_21
cc_57 N_noxref_21_1 N_MM13_g 0.00145084f
cc_58 N_noxref_21_1 N_Y_8 0.0384639f
cc_59 N_noxref_21_1 N_noxref_20_1 0.00177258f
x_PM_AO332x1_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_AO332x1_ASAP7_75t_R%noxref_22
cc_60 N_noxref_22_1 N_NET018_5 0.000511318f
cc_61 N_noxref_22_1 N_NET018_14 0.0374057f
cc_62 N_noxref_22_1 N_MM1_g 0.00145454f
cc_63 N_noxref_22_1 N_NET030_12 0.000471055f
x_PM_AO332x1_ASAP7_75t_R%C2 VSS C2 N_MM0_g N_C2_4 N_C2_1
+ PM_AO332x1_ASAP7_75t_R%C2
cc_64 N_MM0_g N_NET018_5 0.00024254f
cc_65 N_MM0_g N_NET018_4 0.00125312f
cc_66 N_C2_4 N_NET018_20 0.000574623f
cc_67 N_C2_1 N_NET018_15 0.000870849f
cc_68 N_C2_4 N_NET018_19 0.00124633f
cc_69 N_C2_4 N_NET018_4 0.00215805f
cc_70 N_MM0_g N_NET018_15 0.0353316f
cc_71 N_MM0_g N_B3_1 0.000847772f
cc_72 N_C2_4 N_B3_4 0.00324406f
cc_73 N_MM0_g N_MM4_g 0.00402815f
x_PM_AO332x1_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_AO332x1_ASAP7_75t_R%noxref_23
cc_74 N_noxref_23_1 N_NET018_21 0.000237481f
cc_75 N_noxref_23_1 N_NET018_15 0.000988568f
cc_76 N_noxref_23_1 N_MM1_g 0.00143854f
cc_77 N_noxref_23_1 N_NET030_12 0.0359715f
cc_78 N_noxref_23_1 N_noxref_22_1 0.00176902f
x_PM_AO332x1_ASAP7_75t_R%B1 VSS B1 N_MM6_g N_B1_1 N_B1_4
+ PM_AO332x1_ASAP7_75t_R%B1
cc_79 N_B1_1 N_NET018_13 0.000857628f
cc_80 N_B1_4 N_NET018_19 0.00124886f
cc_81 N_MM6_g N_NET018_3 0.00155679f
cc_82 N_B1_4 N_NET018_3 0.00182046f
cc_83 N_MM6_g N_NET018_13 0.0356814f
cc_84 N_B1_1 N_MM9_g 0.000859922f
cc_85 N_B1_4 N_A1_4 0.0030526f
cc_86 N_MM6_g N_MM9_g 0.00401436f
x_PM_AO332x1_ASAP7_75t_R%B3 VSS B3 N_MM4_g N_B3_4 N_B3_1
+ PM_AO332x1_ASAP7_75t_R%B3
cc_87 N_B3_4 N_NET018_19 0.00307354f
cc_88 N_B3_1 N_B2_1 0.00134943f
cc_89 N_B3_4 N_B2_4 0.00334639f
cc_90 N_MM4_g N_MM5_g 0.00613f
x_PM_AO332x1_ASAP7_75t_R%Y VSS Y N_MM13_d N_MM15_d N_Y_7 N_Y_2 N_Y_1 N_Y_8
+ N_Y_10 N_Y_9 PM_AO332x1_ASAP7_75t_R%Y
cc_91 N_Y_7 N_NET018_22 0.00016414f
cc_92 N_Y_7 N_NET018_23 0.000303145f
cc_93 N_Y_7 N_NET018_17 0.000729301f
cc_94 N_Y_7 N_NET018_1 0.000806441f
cc_95 N_Y_2 N_MM13_g 0.00107008f
cc_96 N_Y_1 N_MM13_g 0.00142399f
cc_97 N_Y_8 N_NET018_1 0.00160859f
cc_98 N_Y_10 N_NET018_22 0.00334478f
cc_99 N_Y_9 N_NET018_16 0.0045492f
cc_100 N_Y_8 N_MM13_g 0.0152364f
cc_101 N_Y_7 N_MM13_g 0.0549099f
x_PM_AO332x1_ASAP7_75t_R%C1 VSS C1 N_MM1_g N_C1_1 N_C1_4
+ PM_AO332x1_ASAP7_75t_R%C1
cc_102 N_MM1_g N_NET018_15 0.0157287f
cc_103 N_C1_1 N_NET018_5 0.000895478f
cc_104 N_MM1_g N_NET018_4 0.000944882f
cc_105 N_C1_4 N_NET018_20 0.00109606f
cc_106 N_C1_4 N_NET018_19 0.0011243f
cc_107 N_C1_1 N_NET018_14 0.00167051f
cc_108 N_MM1_g N_NET018_5 0.00167795f
cc_109 N_C1_4 N_NET018_21 0.00666596f
cc_110 N_MM1_g N_NET018_14 0.0546979f
cc_111 N_C1_1 N_C2_1 0.00116073f
cc_112 N_C1_4 N_C2_4 0.00333415f
cc_113 N_MM1_g N_MM0_g 0.00581218f
x_PM_AO332x1_ASAP7_75t_R%A1 VSS A1 N_MM9_g N_A1_1 N_A1_4
+ PM_AO332x1_ASAP7_75t_R%A1
cc_114 N_A1_1 N_NET018_13 0.000869579f
cc_115 N_A1_4 N_NET018_19 0.00124385f
cc_116 N_MM9_g N_NET018_3 0.00155614f
cc_117 N_A1_4 N_NET018_3 0.00178172f
cc_118 N_MM9_g N_NET018_13 0.03571f
cc_119 N_A1_1 N_A2_1 0.00126013f
cc_120 N_A1_4 N_A2_4 0.00364929f
cc_121 N_MM9_g N_MM8_g 0.00619523f
x_PM_AO332x1_ASAP7_75t_R%B2 VSS B2 N_MM5_g N_B2_4 N_B2_1
+ PM_AO332x1_ASAP7_75t_R%B2
cc_122 N_B2_4 N_NET018_3 0.000274794f
cc_123 N_B2_4 N_NET018_13 0.000407238f
cc_124 N_B2_4 N_NET018_19 0.00333653f
cc_125 N_B2_1 N_B1_1 0.0013338f
cc_126 N_B2_4 N_B1_4 0.00338495f
cc_127 N_MM5_g N_MM6_g 0.00598632f
x_PM_AO332x1_ASAP7_75t_R%NET018 VSS N_MM13_g N_MM14_d N_MM12_d N_MM17_d N_MM0_d
+ N_MM1_d N_NET018_17 N_NET018_24 N_NET018_1 N_NET018_16 N_NET018_13
+ N_NET018_18 N_NET018_3 N_NET018_19 N_NET018_5 N_NET018_4 N_NET018_20
+ N_NET018_15 N_NET018_14 N_NET018_21 N_NET018_22 N_NET018_23 N_NET018_26
+ PM_AO332x1_ASAP7_75t_R%NET018
x_PM_AO332x1_ASAP7_75t_R%NET030 VSS N_MM6_d N_MM5_d N_MM4_d N_MM0_s N_MM1_s
+ N_NET030_13 N_NET030_3 N_NET030_12 N_NET030_2 N_NET030_10 N_NET030_1
+ N_NET030_11 PM_AO332x1_ASAP7_75t_R%NET030
cc_128 N_NET030_13 N_NET018_5 0.000133981f
cc_129 N_NET030_13 N_NET018_4 0.00121896f
cc_130 N_NET030_13 N_NET018_15 0.000560771f
cc_131 N_NET030_13 N_NET018_26 0.00064463f
cc_132 N_NET030_3 N_NET018_20 0.000665905f
cc_133 N_NET030_3 N_NET018_21 0.000701942f
cc_134 N_NET030_12 N_NET018_15 0.00188102f
cc_135 N_NET030_2 N_NET018_4 0.0013421f
cc_136 N_NET030_3 N_NET018_4 0.00529195f
cc_137 N_NET030_13 N_NET018_20 0.00816444f
cc_138 N_NET030_10 N_B1_1 0.000580185f
cc_139 N_NET030_1 N_MM6_g 0.000906067f
cc_140 N_NET030_10 N_MM6_g 0.0337731f
cc_141 N_NET030_10 N_B2_1 0.000732578f
cc_142 N_NET030_1 N_MM5_g 0.000910373f
cc_143 N_NET030_10 N_MM5_g 0.0340849f
cc_144 N_NET030_11 N_B3_1 0.000742676f
cc_145 N_NET030_2 N_MM4_g 0.000939576f
cc_146 N_NET030_11 N_MM4_g 0.0343067f
cc_147 N_NET030_11 N_C2_1 0.000728182f
cc_148 N_NET030_2 N_MM0_g 0.000941806f
cc_149 N_NET030_11 N_MM0_g 0.0343744f
cc_150 N_NET030_12 N_C1_1 0.000733047f
cc_151 N_NET030_3 N_MM1_g 0.00100978f
cc_152 N_NET030_12 N_MM1_g 0.0341945f
cc_153 N_NET030_11 N_NET031_15 0.000555318f
cc_154 N_NET030_13 N_NET031_3 0.000748731f
cc_155 N_NET030_1 N_NET031_15 0.00082161f
cc_156 N_NET030_11 N_NET031_12 0.00111425f
cc_157 N_NET030_10 N_NET031_12 0.0011164f
cc_158 N_NET030_1 N_NET031_2 0.00123375f
cc_159 N_NET030_1 N_NET031_3 0.00303939f
cc_160 N_NET030_2 N_NET031_3 0.00411672f
cc_161 N_NET030_13 N_NET031_15 0.0100618f
*END of AO332x1_ASAP7_75t_R.pxi
.ENDS
** Design:	AO332x2_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AO332x2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AO332x2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AO332x2_ASAP7_75t_R%NET25 VSS 2 3 1
c1 1 VSS 0.00100184f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2160 $Y2=0.0675
.ends

.subckt PM_AO332x2_ASAP7_75t_R%NET064 VSS 2 3 1
c1 1 VSS 0.000973808f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4320 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4320 $Y2=0.0675
.ends

.subckt PM_AO332x2_ASAP7_75t_R%NET063 VSS 2 3 1
c1 1 VSS 0.000955248f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3780 $Y2=0.0675
.ends

.subckt PM_AO332x2_ASAP7_75t_R%NET26 VSS 2 3 1
c1 1 VSS 0.000974979f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2700 $Y2=0.0675
.ends

.subckt PM_AO332x2_ASAP7_75t_R%NET061 VSS 2 3 1
c1 1 VSS 0.00102269f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.0675 $X2=0.5400 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.0675 $X2=0.5400 $Y2=0.0675
.ends

.subckt PM_AO332x2_ASAP7_75t_R%A3 VSS 6 3 1 4
c1 1 VSS 0.00785514f
c2 3 VSS 0.0836413f
c3 4 VSS 0.00533348f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1207 $X2=0.1890 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1150 $X2=0.1890 $Y2=0.1207
r3 6 4 1.10765 $w=1.3e-08 $l=4.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1150 $X2=0.1890 $Y2=0.1102
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AO332x2_ASAP7_75t_R%A1 VSS 6 3 1 4
c1 1 VSS 0.00762154f
c2 3 VSS 0.0459511f
c3 4 VSS 0.00410412f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1207 $X2=0.2970 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1150 $X2=0.2970 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1150 $X2=0.2970 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_AO332x2_ASAP7_75t_R%A2 VSS 6 3 4 1
c1 1 VSS 0.00663766f
c2 3 VSS 0.0464883f
c3 4 VSS 0.00496394f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1207 $X2=0.2430 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1150 $X2=0.2430 $Y2=0.1207
r3 6 4 1.10765 $w=1.3e-08 $l=4.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1150 $X2=0.2430 $Y2=0.1102
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AO332x2_ASAP7_75t_R%C1 VSS 6 3 1 4
c1 1 VSS 0.00718454f
c2 3 VSS 0.00878249f
c3 4 VSS 0.00450355f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1207 $X2=0.5670 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1150 $X2=0.5670 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1150 $X2=0.5670 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1350
+ $X2=0.5670 $Y2=0.1350
.ends

.subckt PM_AO332x2_ASAP7_75t_R%B2 VSS 6 3 4 1
c1 1 VSS 0.00734344f
c2 3 VSS 0.00981319f
c3 4 VSS 0.00480315f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1207 $X2=0.4050 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1150 $X2=0.4050 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1150 $X2=0.4050 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
.ends

.subckt PM_AO332x2_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.00477162f
.ends

.subckt PM_AO332x2_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.00609647f
.ends

.subckt PM_AO332x2_ASAP7_75t_R%C2 VSS 6 3 4 1
c1 1 VSS 0.00665235f
c2 3 VSS 0.0462288f
c3 4 VSS 0.00457235f
r1 7 8 3.43955 $w=1.3e-08 $l=1.48e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1202 $X2=0.5130 $Y2=0.1350
r2 6 7 1.45744 $w=1.3e-08 $l=6.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1140 $X2=0.5130 $Y2=0.1202
r3 6 4 5.18847 $w=1.3e-08 $l=2.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1140 $X2=0.5130 $Y2=0.0917
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.1350
+ $X2=0.5130 $Y2=0.1350
.ends

.subckt PM_AO332x2_ASAP7_75t_R%B3 VSS 6 3 4 1
c1 1 VSS 0.00821788f
c2 3 VSS 0.0469151f
c3 4 VSS 0.0052599f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1207 $X2=0.4590 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1150 $X2=0.4590 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1150 $X2=0.4590 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1350
+ $X2=0.4590 $Y2=0.1350
.ends

.subckt PM_AO332x2_ASAP7_75t_R%B1 VSS 6 3 1 4
c1 1 VSS 0.0075616f
c2 3 VSS 0.00906133f
c3 4 VSS 0.00483983f
r1 7 8 3.20636 $w=1.3e-08 $l=1.38e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1212 $X2=0.3510 $Y2=0.1350
r2 6 7 1.22425 $w=1.3e-08 $l=5.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1160 $X2=0.3510 $Y2=0.1212
r3 6 4 5.42166 $w=1.3e-08 $l=2.33e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1160 $X2=0.3510 $Y2=0.0927
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
.ends

.subckt PM_AO332x2_ASAP7_75t_R%NET030 VSS 16 17 32 33 35 13 11 3 12 2 10 1
c1 1 VSS 0.00462828f
c2 2 VSS 0.00460923f
c3 3 VSS 0.00514184f
c4 10 VSS 0.00220322f
c5 11 VSS 0.00221104f
c6 12 VSS 0.00228923f
c7 13 VSS 0.0221129f
r1 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2025 $X2=0.5920 $Y2=0.2025
r2 35 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.2025 $X2=0.5795 $Y2=0.2025
r3 33 31 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r4 2 31 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r5 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4860 $Y2=0.2025
r6 32 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r7 3 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2025
+ $X2=0.5940 $Y2=0.2340
r8 2 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2025
+ $X2=0.4860 $Y2=0.2340
r9 27 28 9.0944 $w=1.3e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.5550
+ $Y=0.2340 $X2=0.5940 $Y2=0.2340
r10 26 27 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5235
+ $Y=0.2340 $X2=0.5550 $Y2=0.2340
r11 25 26 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.2340 $X2=0.5235 $Y2=0.2340
r12 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4995
+ $Y=0.2340 $X2=0.5130 $Y2=0.2340
r13 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.2340 $X2=0.4995 $Y2=0.2340
r14 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4725
+ $Y=0.2340 $X2=0.4860 $Y2=0.2340
r15 21 22 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4725 $Y2=0.2340
r16 20 21 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4485
+ $Y=0.2340 $X2=0.4590 $Y2=0.2340
r17 19 20 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4170
+ $Y=0.2340 $X2=0.4485 $Y2=0.2340
r18 18 19 9.0944 $w=1.3e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.4170 $Y2=0.2340
r19 13 18 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3655
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r20 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.2340
r21 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r22 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r23 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3780 $Y2=0.2025
r24 16 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
.ends

.subckt PM_AO332x2_ASAP7_75t_R%NET031 VSS 20 21 38 39 42 43 10 1 13 11 2 15 12 3
c1 1 VSS 0.00993719f
c2 2 VSS 0.00570224f
c3 3 VSS 0.00308094f
c4 10 VSS 0.0045241f
c5 11 VSS 0.00333831f
c6 12 VSS 0.00213144f
c7 13 VSS 0.00869526f
c8 14 VSS 0.000553894f
c9 15 VSS 0.00185386f
c10 16 VSS 0.000537999f
c11 17 VSS 0.00239791f
r1 43 41 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r2 3 41 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r3 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r4 42 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r5 39 37 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r6 2 37 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r7 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r8 38 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r9 3 34 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.1980
r10 2 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.1980
r11 33 34 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4185
+ $Y=0.1980 $X2=0.4320 $Y2=0.1980
r12 32 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1980 $X2=0.4185 $Y2=0.1980
r13 31 32 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.3790
+ $Y=0.1980 $X2=0.4050 $Y2=0.1980
r14 30 31 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3610
+ $Y=0.1980 $X2=0.3790 $Y2=0.1980
r15 29 30 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1980 $X2=0.3610 $Y2=0.1980
r16 28 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.1980 $X2=0.3510 $Y2=0.1980
r17 27 28 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1980 $X2=0.3375 $Y2=0.1980
r18 15 27 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3105
+ $Y=0.1980 $X2=0.3240 $Y2=0.1980
r19 15 16 1.40651 $w=1.51875e-08 $l=1.45774e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3105 $Y=0.1980 $X2=0.2970 $Y2=0.2035
r20 14 17 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.2160 $X2=0.2970 $Y2=0.2340
r21 14 16 2.45586 $w=1.44e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.2160 $X2=0.2970 $Y2=0.2035
r22 17 25 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.2340 $X2=0.2700 $Y2=0.2340
r23 24 25 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r24 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.2340 $X2=0.2430 $Y2=0.2340
r25 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2295 $Y2=0.2340
r26 13 22 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2035
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r27 1 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.2340
r28 21 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r29 1 19 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r30 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r31 20 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
.ends

.subckt PM_AO332x2_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.04238f
.ends

.subckt PM_AO332x2_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.0423793f
.ends

.subckt PM_AO332x2_ASAP7_75t_R%Y VSS 23 16 17 31 32 7 8 9 1 2 10
c1 1 VSS 0.0100915f
c2 2 VSS 0.0109641f
c3 7 VSS 0.00457281f
c4 8 VSS 0.00456993f
c5 9 VSS 0.00755249f
c6 10 VSS 0.0116446f
c7 11 VSS 0.00933823f
c8 12 VSS 0.00351954f
c9 13 VSS 0.00348702f
r1 32 30 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r2 2 30 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r4 31 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
r5 2 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.2340
r6 11 27 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0675
+ $Y=0.2340 $X2=0.1080 $Y2=0.2340
r7 11 13 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0675 $Y=0.2340 $X2=0.0270 $Y2=0.2340
r8 13 26 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0270 $Y2=0.2125
r9 25 26 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1755 $X2=0.0270 $Y2=0.2125
r10 24 25 6.99569 $w=1.3e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1455 $X2=0.0270 $Y2=0.1755
r11 23 24 1.39914 $w=1.3e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1395 $X2=0.0270 $Y2=0.1455
r12 23 22 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1395 $X2=0.0270 $Y2=0.1010
r13 9 12 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0540 $X2=0.0270 $Y2=0.0360
r14 9 22 10.9599 $w=1.3e-08 $l=4.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0540 $X2=0.0270 $Y2=0.1010
r15 10 18 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0675
+ $Y=0.0360 $X2=0.1080 $Y2=0.0360
r16 10 12 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0675 $Y=0.0360 $X2=0.0270 $Y2=0.0360
r17 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1080 $Y2=0.0360
r18 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r19 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r20 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r21 16 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.0935 $Y2=0.0675
.ends

.subckt PM_AO332x2_ASAP7_75t_R%NET018 VSS 12 13 67 68 72 80 81 18 25 1 17 14 19
+ 3 20 5 4 21 16 22 15 23 24 27
c1 1 VSS 0.00784065f
c2 3 VSS 0.00586999f
c3 4 VSS 0.00284371f
c4 5 VSS 0.00602665f
c5 12 VSS 0.0808061f
c6 13 VSS 0.0806144f
c7 14 VSS 0.00458116f
c8 15 VSS 0.00453825f
c9 16 VSS 0.00389171f
c10 17 VSS 0.00236515f
c11 18 VSS 0.00144118f
c12 19 VSS 0.000687747f
c13 20 VSS 0.0400233f
c14 21 VSS 0.00133154f
c15 22 VSS 0.00510512f
c16 23 VSS 0.000542418f
c17 24 VSS 0.0027649f
c18 25 VSS 0.000657172f
c19 26 VSS 0.00325461f
c20 27 VSS 0.00138553f
r1 81 79 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r2 4 79 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5400 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r3 16 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.2025 $X2=0.5400 $Y2=0.2025
r4 80 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.2025 $X2=0.5255 $Y2=0.2025
r5 4 76 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.2025
+ $X2=0.5400 $Y2=0.1980
r6 76 77 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1980 $X2=0.5535 $Y2=0.1980
r7 74 77 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1980 $X2=0.5535 $Y2=0.1980
r8 73 74 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.5930
+ $Y=0.1980 $X2=0.5670 $Y2=0.1980
r9 21 27 0.682785 $w=1.75e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6110
+ $Y=0.1980 $X2=0.6210 $Y2=0.1980
r10 21 73 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6110
+ $Y=0.1980 $X2=0.5930 $Y2=0.1980
r11 27 70 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.1980 $X2=0.6210 $Y2=0.1765
r12 15 5 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.0675 $X2=0.5920 $Y2=0.0675
r13 72 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0675 $X2=0.5795 $Y2=0.0675
r14 69 70 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1170 $X2=0.6210 $Y2=0.1765
r15 22 26 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.0575 $X2=0.6210 $Y2=0.0360
r16 22 69 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0575 $X2=0.6210 $Y2=0.1170
r17 68 66 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r18 3 66 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r19 14 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3240 $Y2=0.0675
r20 67 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r21 5 63 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0675
+ $X2=0.5940 $Y2=0.0360
r22 26 64 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.0360 $X2=0.6075 $Y2=0.0360
r23 3 49 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0675
+ $X2=0.3240 $Y2=0.0360
r24 63 64 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0360 $X2=0.6075 $Y2=0.0360
r25 62 63 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5805
+ $Y=0.0360 $X2=0.5940 $Y2=0.0360
r26 61 62 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0360 $X2=0.5805 $Y2=0.0360
r27 60 61 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.5415
+ $Y=0.0360 $X2=0.5670 $Y2=0.0360
r28 59 60 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5235
+ $Y=0.0360 $X2=0.5415 $Y2=0.0360
r29 58 59 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0360 $X2=0.5235 $Y2=0.0360
r30 57 58 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.0360 $X2=0.5130 $Y2=0.0360
r31 56 57 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0360 $X2=0.4860 $Y2=0.0360
r32 55 56 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4485
+ $Y=0.0360 $X2=0.4590 $Y2=0.0360
r33 54 55 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4305
+ $Y=0.0360 $X2=0.4485 $Y2=0.0360
r34 53 54 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0360 $X2=0.4305 $Y2=0.0360
r35 52 53 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0360 $X2=0.4050 $Y2=0.0360
r36 51 52 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r37 50 51 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.0360 $X2=0.3510 $Y2=0.0360
r38 49 50 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.0360 $X2=0.3375 $Y2=0.0360
r39 48 49 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3105
+ $Y=0.0360 $X2=0.3240 $Y2=0.0360
r40 47 48 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.3105 $Y2=0.0360
r41 46 47 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.2970 $Y2=0.0360
r42 45 46 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r43 44 45 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2170
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r44 20 24 0.682785 $w=1.75e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1990
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r45 20 44 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1990
+ $Y=0.0360 $X2=0.2170 $Y2=0.0360
r46 19 25 2.45586 $w=1.44e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0540 $X2=0.1890 $Y2=0.0665
r47 19 24 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0540 $X2=0.1890 $Y2=0.0360
r48 25 42 4.08819 $w=1.38974e-08 $l=2.55979e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0665 $X2=0.1640 $Y2=0.0720
r49 18 23 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1460 $Y=0.0720 $X2=0.1350 $Y2=0.0720
r50 18 42 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1460
+ $Y=0.0720 $X2=0.1640 $Y2=0.0720
r51 23 41 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.0720 $X2=0.1350 $Y2=0.0935
r52 17 39 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1160 $X2=0.1350 $Y2=0.1350
r53 17 41 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1160 $X2=0.1350 $Y2=0.0935
r54 13 35 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1350 $Y2=0.1350
r55 35 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
r56 34 35 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1255
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r57 32 34 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1350 $X2=0.1255 $Y2=0.1350
r58 31 32 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1350 $X2=0.1225 $Y2=0.1350
r59 30 31 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1350 $X2=0.1080 $Y2=0.1350
r60 12 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r61 1 29 2.90696 $w=2.1681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0705 $Y2=0.1350
r62 1 30 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1350
r63 12 29 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.0810 $Y=0.1350 $X2=0.0705 $Y2=0.1350
r64 12 30 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1350
.ends


*
.SUBCKT AO332x2_ASAP7_75t_R VSS VDD A3 A2 A1 B1 B2 B3 C2 C1 Y
*
* VSS VSS
* VDD VDD
* A3 A3
* A2 A2
* A1 A1
* B1 B1
* B2 B2
* B3 B3
* C2 C2
* C1 C1
* Y Y
*
*

MM13 N_MM13_d N_MM13_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM13@2 N_MM13@2_d N_MM15@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM8_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM14 N_MM14_d N_MM9_g N_MM14_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM12 N_MM12_d N_MM6_g N_MM12_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 N_MM11_d N_MM5_g N_MM11_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM16 N_MM16_d N_MM0_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM17 N_MM17_d N_MM1_g N_MM17_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM15 N_MM15_d N_MM13_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM15@2 N_MM15@2_d N_MM15@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM8_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM6_g N_MM6_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g N_MM4_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM0_g N_MM0_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AO332x2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AO332x2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AO332x2_ASAP7_75t_R%NET25 VSS N_MM3_d N_MM2_s N_NET25_1
+ PM_AO332x2_ASAP7_75t_R%NET25
cc_1 N_NET25_1 N_MM7_g 0.017362f
cc_2 N_NET25_1 N_MM8_g 0.0173107f
x_PM_AO332x2_ASAP7_75t_R%NET064 VSS N_MM11_s N_MM10_d N_NET064_1
+ PM_AO332x2_ASAP7_75t_R%NET064
cc_3 N_NET064_1 N_MM5_g 0.0174138f
cc_4 N_NET064_1 N_MM4_g 0.0172863f
x_PM_AO332x2_ASAP7_75t_R%NET063 VSS N_MM12_s N_MM11_d N_NET063_1
+ PM_AO332x2_ASAP7_75t_R%NET063
cc_5 N_NET063_1 N_MM6_g 0.017319f
cc_6 N_NET063_1 N_MM5_g 0.017287f
x_PM_AO332x2_ASAP7_75t_R%NET26 VSS N_MM2_d N_MM14_s N_NET26_1
+ PM_AO332x2_ASAP7_75t_R%NET26
cc_7 N_NET26_1 N_MM8_g 0.0173382f
cc_8 N_NET26_1 N_MM9_g 0.0172484f
x_PM_AO332x2_ASAP7_75t_R%NET061 VSS N_MM16_d N_MM17_s N_NET061_1
+ PM_AO332x2_ASAP7_75t_R%NET061
cc_9 N_NET061_1 N_MM0_g 0.0174323f
cc_10 N_NET061_1 N_MM1_g 0.0173457f
x_PM_AO332x2_ASAP7_75t_R%A3 VSS A3 N_MM7_g N_A3_1 N_A3_4
+ PM_AO332x2_ASAP7_75t_R%A3
cc_11 N_MM7_g N_NET018_18 0.000395035f
cc_12 N_MM7_g N_NET018_25 0.000606122f
cc_13 N_A3_1 N_NET018_1 0.00192009f
cc_14 N_A3_4 N_NET018_17 0.00319705f
cc_15 N_MM7_g N_MM15@2_g 0.00380966f
x_PM_AO332x2_ASAP7_75t_R%A1 VSS A1 N_MM9_g N_A1_1 N_A1_4
+ PM_AO332x2_ASAP7_75t_R%A1
cc_16 N_MM9_g N_NET018_3 0.00181078f
cc_17 N_A1_1 N_NET018_14 0.000869617f
cc_18 N_A1_4 N_NET018_20 0.00129316f
cc_19 N_A1_4 N_NET018_3 0.0018179f
cc_20 N_MM9_g N_NET018_14 0.0355309f
cc_21 N_A1_1 N_A2_1 0.0013212f
cc_22 N_A1_4 N_A2_4 0.00368813f
cc_23 N_MM9_g N_MM8_g 0.00600184f
x_PM_AO332x2_ASAP7_75t_R%A2 VSS A2 N_MM8_g N_A2_4 N_A2_1
+ PM_AO332x2_ASAP7_75t_R%A2
cc_24 N_A2_4 N_NET018_14 0.000259299f
cc_25 N_A2_4 N_NET018_19 0.000191671f
cc_26 N_A2_4 N_NET018_3 0.00027294f
cc_27 N_MM8_g N_NET018_14 0.000461888f
cc_28 N_A2_4 N_NET018_20 0.00137626f
cc_29 N_A2_4 N_NET018_25 0.00285332f
cc_30 N_A2_1 N_A3_1 0.0012846f
cc_31 N_A2_4 N_A3_4 0.00376518f
cc_32 N_MM8_g N_MM7_g 0.00606155f
x_PM_AO332x2_ASAP7_75t_R%C1 VSS C1 N_MM1_g N_C1_1 N_C1_4
+ PM_AO332x2_ASAP7_75t_R%C1
cc_33 N_MM1_g N_NET018_16 0.0157086f
cc_34 N_C1_1 N_NET018_5 0.000892474f
cc_35 N_MM1_g N_NET018_4 0.000910517f
cc_36 N_C1_4 N_NET018_21 0.0010625f
cc_37 N_C1_4 N_NET018_20 0.0012046f
cc_38 N_MM1_g N_NET018_5 0.00168483f
cc_39 N_C1_1 N_NET018_16 0.00182279f
cc_40 N_C1_4 N_NET018_22 0.00666368f
cc_41 N_MM1_g N_NET018_15 0.0547601f
cc_42 N_C1_1 N_C2_1 0.00119783f
cc_43 N_C1_4 N_C2_4 0.00328442f
cc_44 N_MM1_g N_MM0_g 0.00585946f
x_PM_AO332x2_ASAP7_75t_R%B2 VSS B2 N_MM5_g N_B2_4 N_B2_1
+ PM_AO332x2_ASAP7_75t_R%B2
cc_45 N_B2_4 N_NET018_3 0.000273528f
cc_46 N_B2_4 N_NET018_14 0.00040742f
cc_47 N_B2_4 N_NET018_20 0.00330004f
cc_48 N_B2_1 N_B1_1 0.00136844f
cc_49 N_B2_4 N_B1_4 0.00349424f
cc_50 N_MM5_g N_MM6_g 0.00606401f
x_PM_AO332x2_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_AO332x2_ASAP7_75t_R%noxref_22
cc_51 N_noxref_22_1 N_NET018_5 0.000506533f
cc_52 N_noxref_22_1 N_NET018_15 0.0375055f
cc_53 N_noxref_22_1 N_MM1_g 0.00146127f
cc_54 N_noxref_22_1 N_NET030_12 0.000469041f
x_PM_AO332x2_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_AO332x2_ASAP7_75t_R%noxref_23
cc_55 N_noxref_23_1 N_NET018_22 0.000239083f
cc_56 N_noxref_23_1 N_NET018_16 0.00098706f
cc_57 N_noxref_23_1 N_MM1_g 0.001448f
cc_58 N_noxref_23_1 N_NET030_12 0.0358971f
cc_59 N_noxref_23_1 N_noxref_22_1 0.00177008f
x_PM_AO332x2_ASAP7_75t_R%C2 VSS C2 N_MM0_g N_C2_4 N_C2_1
+ PM_AO332x2_ASAP7_75t_R%C2
cc_60 N_MM0_g N_NET018_5 0.000244522f
cc_61 N_MM0_g N_NET018_4 0.001261f
cc_62 N_C2_4 N_NET018_21 0.000593841f
cc_63 N_C2_1 N_NET018_16 0.000852303f
cc_64 N_C2_4 N_NET018_20 0.00131821f
cc_65 N_C2_4 N_NET018_4 0.0021358f
cc_66 N_MM0_g N_NET018_16 0.0353654f
cc_67 N_C2_4 N_B3_1 0.000846936f
cc_68 N_MM0_g N_MM4_g 0.00326853f
cc_69 N_C2_4 N_B3_4 0.00423418f
x_PM_AO332x2_ASAP7_75t_R%B3 VSS B3 N_MM4_g N_B3_4 N_B3_1
+ PM_AO332x2_ASAP7_75t_R%B3
cc_70 N_B3_4 N_NET018_20 0.00325945f
cc_71 N_B3_1 N_B2_1 0.00134243f
cc_72 N_B3_4 N_B2_4 0.00332981f
cc_73 N_MM4_g N_MM5_g 0.00596617f
x_PM_AO332x2_ASAP7_75t_R%B1 VSS B1 N_MM6_g N_B1_1 N_B1_4
+ PM_AO332x2_ASAP7_75t_R%B1
cc_74 N_B1_1 N_NET018_14 0.000858553f
cc_75 N_B1_4 N_NET018_20 0.00131618f
cc_76 N_MM6_g N_NET018_3 0.00155349f
cc_77 N_B1_4 N_NET018_3 0.00175032f
cc_78 N_MM6_g N_NET018_14 0.0356176f
cc_79 N_B1_1 N_MM9_g 0.000883159f
cc_80 N_B1_4 N_A1_4 0.00316839f
cc_81 N_MM6_g N_MM9_g 0.00401093f
x_PM_AO332x2_ASAP7_75t_R%NET030 VSS N_MM6_d N_MM5_d N_MM4_d N_MM0_s N_MM1_s
+ N_NET030_13 N_NET030_11 N_NET030_3 N_NET030_12 N_NET030_2 N_NET030_10
+ N_NET030_1 PM_AO332x2_ASAP7_75t_R%NET030
cc_82 N_NET030_13 N_NET018_5 0.00013287f
cc_83 N_NET030_13 N_NET018_4 0.000995987f
cc_84 N_NET030_11 N_NET018_16 0.00168234f
cc_85 N_NET030_13 N_NET018_27 0.000639589f
cc_86 N_NET030_3 N_NET018_22 0.000728273f
cc_87 N_NET030_12 N_NET018_16 0.000766395f
cc_88 N_NET030_3 N_NET018_4 0.00249164f
cc_89 N_NET030_2 N_NET018_4 0.00414131f
cc_90 N_NET030_13 N_NET018_21 0.00914809f
cc_91 N_NET030_10 N_B1_1 0.000578731f
cc_92 N_NET030_1 N_MM6_g 0.000906092f
cc_93 N_NET030_10 N_MM6_g 0.0338637f
cc_94 N_NET030_10 N_B2_1 0.000770854f
cc_95 N_NET030_1 N_MM5_g 0.000907019f
cc_96 N_NET030_10 N_MM5_g 0.0339898f
cc_97 N_NET030_11 N_B3_1 0.000730958f
cc_98 N_NET030_2 N_MM4_g 0.000937776f
cc_99 N_NET030_11 N_MM4_g 0.0343943f
cc_100 N_NET030_11 N_C2_1 0.000739572f
cc_101 N_NET030_2 N_MM0_g 0.000936101f
cc_102 N_NET030_11 N_MM0_g 0.0343037f
cc_103 N_NET030_12 N_C1_1 0.000738912f
cc_104 N_NET030_3 N_MM1_g 0.00100672f
cc_105 N_NET030_12 N_MM1_g 0.0341708f
cc_106 N_NET030_11 N_NET031_15 0.000554512f
cc_107 N_NET030_13 N_NET031_3 0.000749985f
cc_108 N_NET030_1 N_NET031_15 0.000820867f
cc_109 N_NET030_10 N_NET031_12 0.00111391f
cc_110 N_NET030_10 N_NET031_11 0.00111489f
cc_111 N_NET030_2 N_NET031_3 0.00132048f
cc_112 N_NET030_1 N_NET031_3 0.0027696f
cc_113 N_NET030_1 N_NET031_2 0.00426658f
cc_114 N_NET030_13 N_NET031_15 0.0102101f
x_PM_AO332x2_ASAP7_75t_R%NET031 VSS N_MM7_d N_MM8_d N_MM9_d N_MM6_s N_MM5_s
+ N_MM4_s N_NET031_10 N_NET031_1 N_NET031_13 N_NET031_11 N_NET031_2 N_NET031_15
+ N_NET031_12 N_NET031_3 PM_AO332x2_ASAP7_75t_R%NET031
cc_115 N_NET031_10 N_A3_1 0.000777555f
cc_116 N_NET031_1 N_A3_4 0.00107511f
cc_117 N_NET031_1 N_MM7_g 0.00115152f
cc_118 N_NET031_10 N_MM7_g 0.034031f
cc_119 N_NET031_10 N_A2_1 0.000664024f
cc_120 N_NET031_13 N_A2_4 0.00100485f
cc_121 N_NET031_1 N_MM8_g 0.00116276f
cc_122 N_NET031_1 N_A2_4 0.00208979f
cc_123 N_NET031_10 N_MM8_g 0.0340297f
cc_124 N_NET031_11 N_A1_4 0.000459353f
cc_125 N_NET031_11 N_A1_1 0.000815324f
cc_126 N_NET031_2 N_MM9_g 0.000849394f
cc_127 N_NET031_2 N_A1_4 0.00106747f
cc_128 N_NET031_11 N_MM9_g 0.0340603f
cc_129 N_NET031_11 N_B1_1 0.000617059f
cc_130 N_NET031_2 N_MM6_g 0.000838826f
cc_131 N_NET031_15 N_B1_4 0.00113999f
cc_132 N_NET031_2 N_B1_4 0.00129311f
cc_133 N_NET031_11 N_MM6_g 0.033515f
cc_134 N_NET031_12 N_B2_1 0.000778657f
cc_135 N_NET031_3 N_MM5_g 0.000899524f
cc_136 N_NET031_15 N_B2_4 0.00114348f
cc_137 N_NET031_3 N_B2_4 0.0012633f
cc_138 N_NET031_12 N_MM5_g 0.0336697f
cc_139 N_NET031_12 N_B3_4 0.000621907f
cc_140 N_NET031_12 N_B3_1 0.000754665f
cc_141 N_NET031_3 N_B3_4 0.000786161f
cc_142 N_NET031_3 N_MM4_g 0.000895322f
cc_143 N_NET031_12 N_MM4_g 0.0333439f
x_PM_AO332x2_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_AO332x2_ASAP7_75t_R%noxref_21
cc_144 N_noxref_21_1 N_MM13_g 0.00146671f
cc_145 N_noxref_21_1 N_Y_8 0.000843538f
cc_146 N_noxref_21_1 N_noxref_20_1 0.0017768f
x_PM_AO332x2_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_AO332x2_ASAP7_75t_R%noxref_20
cc_147 N_noxref_20_1 N_MM13_g 0.00146907f
cc_148 N_noxref_20_1 N_Y_7 0.000844161f
x_PM_AO332x2_ASAP7_75t_R%Y VSS Y N_MM13_d N_MM13@2_d N_MM15_d N_MM15@2_d N_Y_7
+ N_Y_8 N_Y_9 N_Y_1 N_Y_2 N_Y_10 PM_AO332x2_ASAP7_75t_R%Y
cc_149 N_Y_7 N_NET018_23 0.000231837f
cc_150 N_Y_7 N_NET018_24 0.000248312f
cc_151 N_Y_7 N_NET018_17 0.000284558f
cc_152 N_Y_7 N_NET018_1 0.000464874f
cc_153 N_Y_7 N_NET018_18 0.000697366f
cc_154 N_Y_8 N_MM13_g 0.0309788f
cc_155 N_Y_9 N_NET018_1 0.000929087f
cc_156 N_Y_1 N_NET018_17 0.00141858f
cc_157 N_Y_2 N_MM13_g 0.00195935f
cc_158 N_Y_1 N_MM13_g 0.0023578f
cc_159 N_Y_10 N_NET018_23 0.00329342f
cc_160 N_Y_8 N_NET018_1 0.00476751f
cc_161 N_Y_7 N_MM15@2_g 0.0372187f
cc_162 N_Y_7 N_MM13_g 0.0684942f
x_PM_AO332x2_ASAP7_75t_R%NET018 VSS N_MM13_g N_MM15@2_g N_MM14_d N_MM12_d
+ N_MM17_d N_MM0_d N_MM1_d N_NET018_18 N_NET018_25 N_NET018_1 N_NET018_17
+ N_NET018_14 N_NET018_19 N_NET018_3 N_NET018_20 N_NET018_5 N_NET018_4
+ N_NET018_21 N_NET018_16 N_NET018_22 N_NET018_15 N_NET018_23 N_NET018_24
+ N_NET018_27 PM_AO332x2_ASAP7_75t_R%NET018
*END of AO332x2_ASAP7_75t_R.pxi
.ENDS
** Design:	AO333x1_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AO333x1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AO333x1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AO333x1_ASAP7_75t_R%NET54 VSS 2 3 1
c1 1 VSS 0.000992833f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4860 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0675 $X2=0.4860 $Y2=0.0675
.ends

.subckt PM_AO333x1_ASAP7_75t_R%NET55 VSS 2 3 1
c1 1 VSS 0.000961615f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.0675 $X2=0.5400 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.0675 $X2=0.5400 $Y2=0.0675
.ends

.subckt PM_AO333x1_ASAP7_75t_R%NET58 VSS 2 3 1
c1 1 VSS 0.000982349f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_AO333x1_ASAP7_75t_R%NET57 VSS 2 3 1
c1 1 VSS 0.000989606f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3780 $Y2=0.0675
.ends

.subckt PM_AO333x1_ASAP7_75t_R%NET59 VSS 2 3 1
c1 1 VSS 0.00100742f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2160 $Y2=0.0675
.ends

.subckt PM_AO333x1_ASAP7_75t_R%NET56 VSS 2 3 1
c1 1 VSS 0.000997942f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3240 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3240 $Y2=0.0675
.ends

.subckt PM_AO333x1_ASAP7_75t_R%NET24 VSS 16 17 33 34 37 38 10 1 13 2 11 12 3
c1 1 VSS 0.0100009f
c2 2 VSS 0.0068487f
c3 3 VSS 0.00460356f
c4 10 VSS 0.00452189f
c5 11 VSS 0.00333145f
c6 12 VSS 0.00213119f
c7 13 VSS 0.0220827f
r1 38 36 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r2 3 36 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r3 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3780 $Y2=0.2025
r4 37 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r5 34 32 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r6 2 32 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r7 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r8 33 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r9 3 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.2340
r10 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.2340
r11 28 29 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3395
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r12 27 28 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3080
+ $Y=0.2340 $X2=0.3395 $Y2=0.2340
r13 26 27 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.2340 $X2=0.3080 $Y2=0.2340
r14 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2835
+ $Y=0.2340 $X2=0.2970 $Y2=0.2340
r15 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.2835 $Y2=0.2340
r16 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r17 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2565 $Y2=0.2340
r18 21 22 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2430 $Y2=0.2340
r19 20 21 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r20 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1755
+ $Y=0.2340 $X2=0.1890 $Y2=0.2340
r21 18 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r22 13 18 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1505
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r23 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r24 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r25 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r26 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r27 16 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
.ends

.subckt PM_AO333x1_ASAP7_75t_R%A1 VSS 6 3 4 1
c1 1 VSS 0.00748373f
c2 3 VSS 0.0459882f
c3 4 VSS 0.00541876f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.0980
r2 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AO333x1_ASAP7_75t_R%B2 VSS 8 3 4 1
c1 1 VSS 0.00748324f
c2 3 VSS 0.00989341f
c3 4 VSS 0.00499996f
r1 9 10 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1055 $X2=0.3510 $Y2=0.1350
r2 8 9 4.89699 $w=1.3e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0845 $X2=0.3510 $Y2=0.1055
r3 8 4 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0845 $X2=0.3510 $Y2=0.0770
r4 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r5 1 10 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
.ends

.subckt PM_AO333x1_ASAP7_75t_R%Y VSS 20 14 28 7 2 1 8 10 9
c1 1 VSS 0.0080659f
c2 2 VSS 0.00906217f
c3 7 VSS 0.00386393f
c4 8 VSS 0.00382447f
c5 9 VSS 0.00395965f
c6 10 VSS 0.00440843f
c7 11 VSS 0.00286529f
c8 12 VSS 0.00635727f
r1 28 27 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r2 8 27 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r3 2 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r4 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r5 12 23 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0270 $Y2=0.2125
r6 12 24 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0405 $Y2=0.2340
r7 22 23 8.51143 $w=1.3e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1760 $X2=0.0270 $Y2=0.2125
r8 21 22 6.99569 $w=1.3e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1460 $X2=0.0270 $Y2=0.1760
r9 20 21 1.51573 $w=1.3e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1395 $X2=0.0270 $Y2=0.1460
r10 20 19 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1395 $X2=0.0270 $Y2=0.1010
r11 9 11 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0540 $X2=0.0270 $Y2=0.0360
r12 9 19 10.9599 $w=1.3e-08 $l=4.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0540 $X2=0.0270 $Y2=0.1010
r13 10 15 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r14 10 11 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0405 $Y=0.0360 $X2=0.0270 $Y2=0.0360
r15 1 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0540 $Y2=0.0360
r16 14 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r17 7 13 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r18 2 8 1e-05
r19 1 7 1e-05
.ends

.subckt PM_AO333x1_ASAP7_75t_R%A3 VSS 8 3 1 4
c1 1 VSS 0.00825553f
c2 3 VSS 0.0838048f
c3 4 VSS 0.00557522f
r1 8 7 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1485 $X2=0.1350 $Y2=0.1460
r2 6 7 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1460
r3 4 6 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1160 $X2=0.1350 $Y2=0.1350
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r5 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AO333x1_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.00476571f
.ends

.subckt PM_AO333x1_ASAP7_75t_R%C3 VSS 8 3 4 1
c1 1 VSS 0.00789942f
c2 3 VSS 0.0467601f
c3 4 VSS 0.00506745f
r1 9 10 6.99569 $w=1.3e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1050 $X2=0.4590 $Y2=0.1350
r2 8 9 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0835 $X2=0.4590 $Y2=0.1050
r3 8 4 1.63233 $w=1.3e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0835 $X2=0.4590 $Y2=0.0765
r4 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r5 1 10 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1350
+ $X2=0.4590 $Y2=0.1350
.ends

.subckt PM_AO333x1_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.00466302f
.ends

.subckt PM_AO333x1_ASAP7_75t_R%B3 VSS 8 3 1 4
c1 1 VSS 0.00796477f
c2 3 VSS 0.00926092f
c3 4 VSS 0.00504261f
r1 8 7 1.28254 $w=1.3e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1545 $X2=0.2970 $Y2=0.1490
r2 6 7 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1490
r3 4 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0980 $X2=0.2970 $Y2=0.1350
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r5 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_AO333x1_ASAP7_75t_R%A2 VSS 10 3 4 1
c1 1 VSS 0.00662097f
c2 3 VSS 0.0463699f
c3 4 VSS 0.0047488f
r1 10 9 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1865 $X2=0.1890 $Y2=0.1650
r2 8 9 6.99569 $w=1.3e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1650
r3 7 8 4.4306 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1160 $X2=0.1890 $Y2=0.1350
r4 4 7 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0935 $X2=0.1890 $Y2=0.1160
r5 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r6 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AO333x1_ASAP7_75t_R%B1 VSS 10 3 4 1
c1 1 VSS 0.00798774f
c2 3 VSS 0.0468235f
c3 4 VSS 0.00509035f
r1 10 9 1.39914 $w=1.3e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1555 $X2=0.4050 $Y2=0.1495
r2 8 9 3.38125 $w=1.3e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1495
r3 4 8 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0980 $X2=0.4050 $Y2=0.1350
r4 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
.ends

.subckt PM_AO333x1_ASAP7_75t_R%C1 VSS 8 3 1 4
c1 1 VSS 0.00689362f
c2 3 VSS 0.00848272f
c3 4 VSS 0.00415793f
r1 9 10 7.22888 $w=1.3e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1040 $X2=0.5670 $Y2=0.1350
r2 8 9 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0815 $X2=0.5670 $Y2=0.1040
r3 8 4 1.39914 $w=1.3e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0815 $X2=0.5670 $Y2=0.0755
r4 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1350
r5 1 10 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1350
+ $X2=0.5670 $Y2=0.1350
.ends

.subckt PM_AO333x1_ASAP7_75t_R%C2 VSS 10 3 1 4
c1 1 VSS 0.0063637f
c2 3 VSS 0.00931693f
c3 4 VSS 0.0041461f
r1 10 9 1.16595 $w=1.3e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1535 $X2=0.5130 $Y2=0.1485
r2 8 9 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1485
r3 4 8 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0980 $X2=0.5130 $Y2=0.1350
r4 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.1350
+ $X2=0.5130 $Y2=0.1350
.ends

.subckt PM_AO333x1_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.00490904f
.ends

.subckt PM_AO333x1_ASAP7_75t_R%NET22 VSS 16 17 37 38 41 42 13 12 3 2 10 1 11
c1 1 VSS 0.00277104f
c2 2 VSS 0.00318144f
c3 3 VSS 0.00274412f
c4 10 VSS 0.00212282f
c5 11 VSS 0.00210812f
c6 12 VSS 0.00209822f
c7 13 VSS 0.00318398f
r1 42 40 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r2 3 40 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5400 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r3 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.2025 $X2=0.5400 $Y2=0.2025
r4 41 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.2025 $X2=0.5255 $Y2=0.2025
r5 38 36 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r6 2 36 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r7 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r8 37 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r9 3 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.2025
+ $X2=0.5400 $Y2=0.1980
r10 2 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.1980
r11 31 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5265
+ $Y=0.1980 $X2=0.5400 $Y2=0.1980
r12 30 31 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1980 $X2=0.5265 $Y2=0.1980
r13 29 30 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.4875
+ $Y=0.1980 $X2=0.5130 $Y2=0.1980
r14 28 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4695
+ $Y=0.1980 $X2=0.4875 $Y2=0.1980
r15 27 28 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1980 $X2=0.4695 $Y2=0.1980
r16 26 27 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4455
+ $Y=0.1980 $X2=0.4590 $Y2=0.1980
r17 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.1980 $X2=0.4455 $Y2=0.1980
r18 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4185
+ $Y=0.1980 $X2=0.4320 $Y2=0.1980
r19 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1980 $X2=0.4185 $Y2=0.1980
r20 22 23 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3955
+ $Y=0.1980 $X2=0.4050 $Y2=0.1980
r21 21 22 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3775
+ $Y=0.1980 $X2=0.3955 $Y2=0.1980
r22 20 21 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1980 $X2=0.3775 $Y2=0.1980
r23 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.1980 $X2=0.3510 $Y2=0.1980
r24 18 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1980 $X2=0.3375 $Y2=0.1980
r25 13 18 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3125
+ $Y=0.1980 $X2=0.3240 $Y2=0.1980
r26 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.1980
r27 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r28 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r29 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r30 16 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
.ends

.subckt PM_AO333x1_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.00453853f
.ends

.subckt PM_AO333x1_ASAP7_75t_R%NET40 VSS 15 60 61 67 74 77 78 21 28 1 20 16 22
+ 3 23 4 18 25 5 19 6 17 27 26 24
c1 1 VSS 0.00351953f
c2 3 VSS 0.00586572f
c3 4 VSS 0.00474009f
c4 5 VSS 0.00563853f
c5 6 VSS 0.00528123f
c6 15 VSS 0.0800143f
c7 16 VSS 0.00300533f
c8 17 VSS 0.00279421f
c9 18 VSS 0.00227996f
c10 19 VSS 0.00242106f
c11 20 VSS 0.00140524f
c12 21 VSS 0.00136994f
c13 22 VSS 0.000665037f
c14 23 VSS 0.0428572f
c15 24 VSS 0.0120399f
c16 25 VSS 0.00297424f
c17 26 VSS 0.000512968f
c18 27 VSS 0.00296012f
c19 28 VSS 0.000665918f
c20 29 VSS 0.00282359f
c21 30 VSS 0.0028693f
r1 78 76 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r2 4 76 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r3 18 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4860 $Y2=0.2025
r4 77 18 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r5 19 6 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2025 $X2=0.5920 $Y2=0.2025
r6 74 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.2025 $X2=0.5795 $Y2=0.2025
r7 4 71 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2025
+ $X2=0.4860 $Y2=0.2340
r8 6 68 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2025
+ $X2=0.5940 $Y2=0.2340
r9 71 72 11.5429 $w=1.3e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.2340 $X2=0.5355 $Y2=0.2340
r10 68 69 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.2340 $X2=0.6075 $Y2=0.2340
r11 24 68 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5805
+ $Y=0.2340 $X2=0.5940 $Y2=0.2340
r12 24 72 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.5805
+ $Y=0.2340 $X2=0.5355 $Y2=0.2340
r13 30 65 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.2340 $X2=0.6210 $Y2=0.2160
r14 30 69 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.2340 $X2=0.6075 $Y2=0.2340
r15 17 5 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.0675 $X2=0.5920 $Y2=0.0675
r16 67 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0675 $X2=0.5795 $Y2=0.0675
r17 64 65 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1980 $X2=0.6210 $Y2=0.2160
r18 63 64 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1765 $X2=0.6210 $Y2=0.1980
r19 62 63 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1170 $X2=0.6210 $Y2=0.1765
r20 25 29 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.0575 $X2=0.6210 $Y2=0.0360
r21 25 62 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0575 $X2=0.6210 $Y2=0.1170
r22 61 59 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r23 3 59 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r24 16 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r25 60 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
r26 5 56 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0675
+ $X2=0.5940 $Y2=0.0360
r27 29 57 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.0360 $X2=0.6075 $Y2=0.0360
r28 3 41 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2700 $Y2=0.0360
r29 56 57 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0360 $X2=0.6075 $Y2=0.0360
r30 55 56 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5805
+ $Y=0.0360 $X2=0.5940 $Y2=0.0360
r31 54 55 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0360 $X2=0.5805 $Y2=0.0360
r32 53 54 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.0360 $X2=0.5670 $Y2=0.0360
r33 52 53 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0360 $X2=0.5400 $Y2=0.0360
r34 51 52 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.0360 $X2=0.5130 $Y2=0.0360
r35 50 51 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0360 $X2=0.4860 $Y2=0.0360
r36 49 50 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4590 $Y2=0.0360
r37 48 49 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r38 47 48 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0360 $X2=0.4050 $Y2=0.0360
r39 46 47 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r40 45 46 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3260
+ $Y=0.0360 $X2=0.3510 $Y2=0.0360
r41 44 45 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3080
+ $Y=0.0360 $X2=0.3260 $Y2=0.0360
r42 43 44 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.3080 $Y2=0.0360
r43 42 43 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2835
+ $Y=0.0360 $X2=0.2970 $Y2=0.0360
r44 41 42 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.2835 $Y2=0.0360
r45 40 41 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r46 39 40 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2565 $Y2=0.0360
r47 38 39 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r48 37 38 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r49 36 37 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1640
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r50 23 27 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1460 $Y=0.0360 $X2=0.1350 $Y2=0.0360
r51 23 36 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1460
+ $Y=0.0360 $X2=0.1640 $Y2=0.0360
r52 22 28 2.45586 $w=1.44e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.0540 $X2=0.1350 $Y2=0.0665
r53 22 27 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0540 $X2=0.1350 $Y2=0.0360
r54 21 26 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0720 $X2=0.0810 $Y2=0.0720
r55 21 28 4.55457 $w=1.3814e-08 $l=2.75545e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0720 $X2=0.1350 $Y2=0.0665
r56 26 34 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0720 $X2=0.0810 $Y2=0.0935
r57 20 32 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1160 $X2=0.0810 $Y2=0.1350
r58 20 34 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1160 $X2=0.0810 $Y2=0.0935
r59 15 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r60 1 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends


*
.SUBCKT AO333x1_ASAP7_75t_R VSS VDD A3 A2 A1 B3 B2 B1 C3 C2 C1 Y
*
* VSS VSS
* VDD VDD
* A3 A3
* A2 A2
* A1 A1
* B3 B3
* B2 B2
* B1 B1
* C3 C3
* C2 C2
* C1 C1
* Y Y
*
*

MM3 N_MM3_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM19 N_MM19_d N_MM17_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM18 N_MM18_d N_MM16_g N_MM18_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM14 N_MM14_d N_MM15_g N_MM14_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM13_g N_MM10_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM12_g N_MM9_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM5_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM6_g N_MM1_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM7_g N_MM0_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM17 N_MM17_d N_MM17_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM16 N_MM16_d N_MM16_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM15 N_MM15_d N_MM15_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM13 N_MM13_d N_MM13_g N_MM13_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM12 N_MM12_d N_MM12_g N_MM12_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 N_MM11_d N_MM11_g N_MM11_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM6_g N_MM6_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM7_g N_MM7_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AO333x1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AO333x1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AO333x1_ASAP7_75t_R%NET54 VSS N_MM2_d N_MM1_s N_NET54_1
+ PM_AO333x1_ASAP7_75t_R%NET54
cc_1 N_NET54_1 N_MM5_g 0.0172749f
cc_2 N_NET54_1 N_MM6_g 0.0174219f
x_PM_AO333x1_ASAP7_75t_R%NET55 VSS N_MM1_d N_MM0_s N_NET55_1
+ PM_AO333x1_ASAP7_75t_R%NET55
cc_3 N_NET55_1 N_MM6_g 0.0173402f
cc_4 N_NET55_1 N_MM7_g 0.0173948f
x_PM_AO333x1_ASAP7_75t_R%NET58 VSS N_MM19_d N_MM18_s N_NET58_1
+ PM_AO333x1_ASAP7_75t_R%NET58
cc_5 N_NET58_1 N_MM17_g 0.0172897f
cc_6 N_NET58_1 N_MM16_g 0.0174157f
x_PM_AO333x1_ASAP7_75t_R%NET57 VSS N_MM9_s N_MM8_d N_NET57_1
+ PM_AO333x1_ASAP7_75t_R%NET57
cc_7 N_NET57_1 N_MM12_g 0.0172975f
cc_8 N_NET57_1 N_MM11_g 0.0174005f
x_PM_AO333x1_ASAP7_75t_R%NET59 VSS N_MM18_d N_MM14_s N_NET59_1
+ PM_AO333x1_ASAP7_75t_R%NET59
cc_9 N_NET59_1 N_MM16_g 0.0172887f
cc_10 N_NET59_1 N_MM15_g 0.0173937f
x_PM_AO333x1_ASAP7_75t_R%NET56 VSS N_MM10_s N_MM9_d N_NET56_1
+ PM_AO333x1_ASAP7_75t_R%NET56
cc_11 N_NET56_1 N_MM13_g 0.0173021f
cc_12 N_NET56_1 N_MM12_g 0.0173881f
x_PM_AO333x1_ASAP7_75t_R%NET24 VSS N_MM17_d N_MM16_d N_MM15_d N_MM13_s N_MM12_s
+ N_MM11_s N_NET24_10 N_NET24_1 N_NET24_13 N_NET24_2 N_NET24_11 N_NET24_12
+ N_NET24_3 PM_AO333x1_ASAP7_75t_R%NET24
cc_13 N_NET24_10 N_A3_1 0.000803875f
cc_14 N_NET24_1 N_A3_4 0.00107688f
cc_15 N_NET24_1 N_MM17_g 0.00117949f
cc_16 N_NET24_10 N_MM17_g 0.0339842f
cc_17 N_NET24_10 N_A2_1 0.000763325f
cc_18 N_NET24_13 N_A2_4 0.00114897f
cc_19 N_NET24_1 N_MM16_g 0.00116557f
cc_20 N_NET24_1 N_A2_4 0.00154513f
cc_21 N_NET24_10 N_MM16_g 0.0335423f
cc_22 N_NET24_2 N_MM15_g 0.00116702f
cc_23 N_NET24_13 N_A1_4 0.00122818f
cc_24 N_NET24_2 N_A1_4 0.00168115f
cc_25 N_NET24_11 N_MM15_g 0.0341602f
cc_26 N_NET24_11 N_B3_1 0.00072029f
cc_27 N_NET24_2 N_MM13_g 0.000922904f
cc_28 N_NET24_11 N_MM13_g 0.033999f
cc_29 N_NET24_12 N_B2_1 0.000654413f
cc_30 N_NET24_3 N_MM12_g 0.000911193f
cc_31 N_NET24_12 N_MM12_g 0.0336296f
cc_32 N_NET24_12 N_B1_1 0.000648938f
cc_33 N_NET24_3 N_MM11_g 0.000900343f
cc_34 N_NET24_12 N_MM11_g 0.0335426f
x_PM_AO333x1_ASAP7_75t_R%A1 VSS A1 N_MM15_g N_A1_4 N_A1_1
+ PM_AO333x1_ASAP7_75t_R%A1
cc_35 N_MM15_g N_NET40_3 0.00183046f
cc_36 N_A1_4 N_NET40_23 0.00120245f
cc_37 N_A1_4 N_NET40_3 0.0018621f
cc_38 N_MM15_g N_NET40_16 0.0362616f
cc_39 N_A1_1 N_A2_1 0.00132093f
cc_40 N_A1_4 N_A2_4 0.00460433f
cc_41 N_MM15_g N_MM16_g 0.0060947f
x_PM_AO333x1_ASAP7_75t_R%B2 VSS B2 N_MM12_g N_B2_4 N_B2_1
+ PM_AO333x1_ASAP7_75t_R%B2
cc_42 N_B2_4 N_NET40_3 0.00027157f
cc_43 N_B2_4 N_NET40_16 0.000401238f
cc_44 N_B2_4 N_NET40_23 0.00333939f
cc_45 N_B2_1 N_B3_1 0.00129781f
cc_46 N_B2_4 N_B3_4 0.00365479f
cc_47 N_MM12_g N_MM13_g 0.00596539f
x_PM_AO333x1_ASAP7_75t_R%Y VSS Y N_MM3_d N_MM4_d N_Y_7 N_Y_2 N_Y_1 N_Y_8 N_Y_10
+ N_Y_9 PM_AO333x1_ASAP7_75t_R%Y
cc_48 N_Y_7 N_NET40_20 0.000130166f
cc_49 N_Y_7 N_NET40_27 0.000155393f
cc_50 N_Y_7 N_NET40_26 0.000223651f
cc_51 N_Y_7 N_NET40_21 0.000396818f
cc_52 N_Y_7 N_NET40_1 0.000768259f
cc_53 N_Y_2 N_MM3_g 0.00108233f
cc_54 N_Y_1 N_MM3_g 0.00143977f
cc_55 N_Y_8 N_NET40_1 0.00160889f
cc_56 N_Y_10 N_NET40_26 0.00265857f
cc_57 N_Y_9 N_NET40_20 0.00462223f
cc_58 N_Y_8 N_MM3_g 0.0154148f
cc_59 N_Y_7 N_MM3_g 0.0545397f
x_PM_AO333x1_ASAP7_75t_R%A3 VSS A3 N_MM17_g N_A3_1 N_A3_4
+ PM_AO333x1_ASAP7_75t_R%A3
cc_60 N_MM17_g N_NET40_21 0.000362774f
cc_61 N_MM17_g N_NET40_28 0.000548258f
cc_62 N_MM17_g N_NET40_1 0.000908257f
cc_63 N_A3_1 N_NET40_1 0.00104873f
cc_64 N_A3_4 N_NET40_20 0.00335344f
cc_65 N_MM17_g N_MM3_g 0.00375143f
x_PM_AO333x1_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_AO333x1_ASAP7_75t_R%noxref_22
cc_66 N_noxref_22_1 N_MM3_g 0.0014586f
cc_67 N_noxref_22_1 N_Y_7 0.0384559f
x_PM_AO333x1_ASAP7_75t_R%C3 VSS C3 N_MM5_g N_C3_4 N_C3_1
+ PM_AO333x1_ASAP7_75t_R%C3
cc_68 N_MM5_g N_NET40_4 0.000928615f
cc_69 N_C3_4 N_NET40_23 0.00126447f
cc_70 N_C3_4 N_NET40_4 0.00164553f
cc_71 N_MM5_g N_NET40_18 0.0356668f
cc_72 N_C3_1 N_B1_1 0.000883509f
cc_73 N_MM5_g N_MM11_g 0.00326679f
cc_74 N_C3_4 N_B1_4 0.00430265f
x_PM_AO333x1_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_AO333x1_ASAP7_75t_R%noxref_23
cc_75 N_noxref_23_1 N_MM3_g 0.00146858f
cc_76 N_noxref_23_1 N_Y_8 0.0385579f
cc_77 N_noxref_23_1 N_noxref_22_1 0.00177186f
x_PM_AO333x1_ASAP7_75t_R%B3 VSS B3 N_MM13_g N_B3_1 N_B3_4
+ PM_AO333x1_ASAP7_75t_R%B3
cc_78 N_MM13_g N_NET40_3 0.00179803f
cc_79 N_B3_1 N_NET40_16 0.000789494f
cc_80 N_B3_4 N_NET40_23 0.0012433f
cc_81 N_B3_4 N_NET40_3 0.00184134f
cc_82 N_MM13_g N_NET40_16 0.0355038f
cc_83 N_B3_1 N_A1_4 0.000886161f
cc_84 N_MM13_g N_MM15_g 0.00327934f
cc_85 N_B3_4 N_A1_4 0.00437769f
x_PM_AO333x1_ASAP7_75t_R%A2 VSS A2 N_MM16_g N_A2_4 N_A2_1
+ PM_AO333x1_ASAP7_75t_R%A2
cc_86 N_A2_4 N_NET40_16 0.000253492f
cc_87 N_A2_4 N_NET40_22 0.000136332f
cc_88 N_A2_4 N_NET40_3 0.000269691f
cc_89 N_MM16_g N_NET40_16 0.000456949f
cc_90 N_A2_4 N_NET40_23 0.0012766f
cc_91 N_A2_4 N_NET40_28 0.00282634f
cc_92 N_A2_1 N_A3_1 0.00136889f
cc_93 N_A2_4 N_A3_4 0.0039372f
cc_94 N_MM16_g N_MM17_g 0.00608168f
x_PM_AO333x1_ASAP7_75t_R%B1 VSS B1 N_MM11_g N_B1_4 N_B1_1
+ PM_AO333x1_ASAP7_75t_R%B1
cc_95 N_B1_4 N_NET40_23 0.0028158f
cc_96 N_B1_1 N_B2_1 0.00125621f
cc_97 N_B1_4 N_B2_4 0.00346126f
cc_98 N_MM11_g N_MM12_g 0.0060244f
x_PM_AO333x1_ASAP7_75t_R%C1 VSS C1 N_MM7_g N_C1_1 N_C1_4
+ PM_AO333x1_ASAP7_75t_R%C1
cc_99 N_MM7_g N_NET40_5 0.00187817f
cc_100 N_MM7_g N_NET40_19 0.015895f
cc_101 N_C1_1 N_NET40_6 0.000836263f
cc_102 N_MM7_g N_NET40_6 0.00108258f
cc_103 N_C1_4 N_NET40_23 0.0011306f
cc_104 N_C1_1 N_NET40_19 0.00169372f
cc_105 N_C1_4 N_NET40_25 0.00614912f
cc_106 N_MM7_g N_NET40_17 0.0546194f
cc_107 N_C1_1 N_C2_1 0.00123918f
cc_108 N_C1_4 N_C2_4 0.00339879f
cc_109 N_MM7_g N_MM6_g 0.00596513f
x_PM_AO333x1_ASAP7_75t_R%C2 VSS C2 N_MM6_g N_C2_1 N_C2_4
+ PM_AO333x1_ASAP7_75t_R%C2
cc_110 N_MM6_g N_NET40_25 0.000121386f
cc_111 N_MM6_g N_NET40_5 0.00027239f
cc_112 N_MM6_g N_NET40_4 0.00122373f
cc_113 N_C2_1 N_NET40_18 0.000815199f
cc_114 N_C2_4 N_NET40_23 0.00139109f
cc_115 N_C2_4 N_NET40_4 0.00162901f
cc_116 N_MM6_g N_NET40_18 0.0353388f
cc_117 N_C2_1 N_C3_1 0.001331f
cc_118 N_C2_4 N_C3_4 0.00350085f
cc_119 N_MM6_g N_MM5_g 0.00600605f
x_PM_AO333x1_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_AO333x1_ASAP7_75t_R%noxref_24
cc_120 N_noxref_24_1 N_NET40_25 0.000320258f
cc_121 N_noxref_24_1 N_NET40_5 0.000504554f
cc_122 N_noxref_24_1 N_NET40_17 0.0375466f
cc_123 N_noxref_24_1 N_MM7_g 0.00145657f
x_PM_AO333x1_ASAP7_75t_R%NET22 VSS N_MM13_d N_MM12_d N_MM11_d N_MM5_s N_MM6_s
+ N_MM7_s N_NET22_13 N_NET22_12 N_NET22_3 N_NET22_2 N_NET22_10 N_NET22_1
+ N_NET22_11 PM_AO333x1_ASAP7_75t_R%NET22
cc_124 N_NET22_13 N_NET40_19 9.75836e-20
cc_125 N_NET22_13 N_NET40_4 0.00112233f
cc_126 N_NET22_13 N_NET40_6 0.000298989f
cc_127 N_NET22_13 N_NET40_18 0.000555089f
cc_128 N_NET22_12 N_NET40_19 0.00167282f
cc_129 N_NET22_13 N_NET40_25 0.000650478f
cc_130 N_NET22_3 N_NET40_24 0.000663094f
cc_131 N_NET22_12 N_NET40_18 0.00111514f
cc_132 N_NET22_2 N_NET40_4 0.00123983f
cc_133 N_NET22_3 N_NET40_4 0.00304636f
cc_134 N_NET22_3 N_NET40_6 0.0042338f
cc_135 N_NET22_13 N_NET40_24 0.0107636f
cc_136 N_NET22_10 N_B3_1 0.000723158f
cc_137 N_NET22_1 N_B3_4 0.000740765f
cc_138 N_NET22_1 N_MM13_g 0.000901424f
cc_139 N_NET22_10 N_MM13_g 0.0339152f
cc_140 N_NET22_10 N_B2_1 0.000702689f
cc_141 N_NET22_1 N_MM12_g 0.000882824f
cc_142 N_NET22_13 N_B2_4 0.0011303f
cc_143 N_NET22_1 N_B2_4 0.00128514f
cc_144 N_NET22_10 N_MM12_g 0.033588f
cc_145 N_NET22_11 N_B1_1 0.000674817f
cc_146 N_NET22_2 N_MM11_g 0.000875373f
cc_147 N_NET22_13 N_B1_4 0.00117565f
cc_148 N_NET22_2 N_B1_4 0.00124483f
cc_149 N_NET22_11 N_MM11_g 0.0335304f
cc_150 N_NET22_2 N_MM5_g 0.000877818f
cc_151 N_NET22_13 N_C3_4 0.00119992f
cc_152 N_NET22_2 N_C3_4 0.00135753f
cc_153 N_NET22_11 N_MM5_g 0.0342648f
cc_154 N_NET22_12 N_C2_1 0.000699073f
cc_155 N_NET22_3 N_MM6_g 0.000862435f
cc_156 N_NET22_13 N_C2_4 0.00116107f
cc_157 N_NET22_3 N_C2_4 0.0012143f
cc_158 N_NET22_12 N_MM6_g 0.0336147f
cc_159 N_NET22_12 N_C1_1 0.000697379f
cc_160 N_NET22_13 N_C1_4 0.000871565f
cc_161 N_NET22_3 N_MM7_g 0.000892569f
cc_162 N_NET22_3 N_C1_4 0.000962123f
cc_163 N_NET22_12 N_MM7_g 0.0335083f
cc_164 N_NET22_10 N_NET24_13 0.000554865f
cc_165 N_NET22_13 N_NET24_3 0.000628031f
cc_166 N_NET22_1 N_NET24_13 0.000775616f
cc_167 N_NET22_10 N_NET24_12 0.00111168f
cc_168 N_NET22_11 N_NET24_12 0.00112031f
cc_169 N_NET22_1 N_NET24_2 0.00133051f
cc_170 N_NET22_1 N_NET24_3 0.00277393f
cc_171 N_NET22_2 N_NET24_3 0.00427909f
cc_172 N_NET22_13 N_NET24_13 0.0105635f
x_PM_AO333x1_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_AO333x1_ASAP7_75t_R%noxref_25
cc_173 N_noxref_25_1 N_NET40_25 0.000319458f
cc_174 N_noxref_25_1 N_NET40_6 0.00050699f
cc_175 N_noxref_25_1 N_NET40_19 0.037758f
cc_176 N_noxref_25_1 N_MM7_g 0.00146163f
cc_177 N_noxref_25_1 N_noxref_24_1 0.0017683f
x_PM_AO333x1_ASAP7_75t_R%NET40 VSS N_MM3_g N_MM14_d N_MM10_d N_MM0_d N_MM7_d
+ N_MM5_d N_MM6_d N_NET40_21 N_NET40_28 N_NET40_1 N_NET40_20 N_NET40_16
+ N_NET40_22 N_NET40_3 N_NET40_23 N_NET40_4 N_NET40_18 N_NET40_25 N_NET40_5
+ N_NET40_19 N_NET40_6 N_NET40_17 N_NET40_27 N_NET40_26 N_NET40_24
+ PM_AO333x1_ASAP7_75t_R%NET40
*END of AO333x1_ASAP7_75t_R.pxi
.ENDS
** Design:	AO333x2_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AO333x2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AO333x2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AO333x2_ASAP7_75t_R%NET54 VSS 2 3 1
c1 1 VSS 0.000991698f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.0675 $X2=0.5400 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.0675 $X2=0.5400 $Y2=0.0675
.ends

.subckt PM_AO333x2_ASAP7_75t_R%NET55 VSS 2 3 1
c1 1 VSS 0.000975057f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.0675 $X2=0.5940 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0675 $X2=0.5940 $Y2=0.0675
.ends

.subckt PM_AO333x2_ASAP7_75t_R%NET59 VSS 2 3 1
c1 1 VSS 0.000993034f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2700 $Y2=0.0675
.ends

.subckt PM_AO333x2_ASAP7_75t_R%NET57 VSS 2 3 1
c1 1 VSS 0.000975584f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4320 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4320 $Y2=0.0675
.ends

.subckt PM_AO333x2_ASAP7_75t_R%NET56 VSS 2 3 1
c1 1 VSS 0.0010072f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3780 $Y2=0.0675
.ends

.subckt PM_AO333x2_ASAP7_75t_R%NET58 VSS 2 3 1
c1 1 VSS 0.000989122f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2160 $Y2=0.0675
.ends

.subckt PM_AO333x2_ASAP7_75t_R%NET24 VSS 16 17 33 34 37 38 1 10 13 2 11 12 3
c1 1 VSS 0.0100723f
c2 2 VSS 0.00696723f
c3 3 VSS 0.00470286f
c4 10 VSS 0.00450949f
c5 11 VSS 0.00332887f
c6 12 VSS 0.00212348f
c7 13 VSS 0.0229118f
r1 38 36 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r2 3 36 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r3 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r4 37 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r5 34 32 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r6 2 32 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r7 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r8 33 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r9 3 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.2340
r10 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.2340
r11 28 29 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3935
+ $Y=0.2340 $X2=0.4320 $Y2=0.2340
r12 27 28 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3620
+ $Y=0.2340 $X2=0.3935 $Y2=0.2340
r13 26 27 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.2340 $X2=0.3620 $Y2=0.2340
r14 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.2340 $X2=0.3510 $Y2=0.2340
r15 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.2340 $X2=0.3375 $Y2=0.2340
r16 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3105
+ $Y=0.2340 $X2=0.3240 $Y2=0.2340
r17 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.2340 $X2=0.3105 $Y2=0.2340
r18 21 22 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.2970 $Y2=0.2340
r19 20 21 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r20 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.2340 $X2=0.2430 $Y2=0.2340
r21 18 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2295 $Y2=0.2340
r22 13 18 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2045
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r23 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.2340
r24 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r25 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r26 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r27 16 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
.ends

.subckt PM_AO333x2_ASAP7_75t_R%A3 VSS 6 3 4 1
c1 1 VSS 0.00803517f
c2 3 VSS 0.0836954f
c3 4 VSS 0.00628494f
r1 7 8 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1095 $X2=0.1890 $Y2=0.1350
r2 6 7 3.96423 $w=1.3e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0925 $X2=0.1890 $Y2=0.1095
r3 6 4 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0925 $X2=0.1890 $Y2=0.0810
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AO333x2_ASAP7_75t_R%A1 VSS 6 3 1 4
c1 1 VSS 0.00753167f
c2 3 VSS 0.0459872f
c3 4 VSS 0.00550511f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.0980
r2 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_AO333x2_ASAP7_75t_R%B3 VSS 8 3 1 4
c1 1 VSS 0.00818228f
c2 3 VSS 0.00938361f
c3 4 VSS 0.00517877f
r1 8 7 1.28254 $w=1.3e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1545 $X2=0.3510 $Y2=0.1490
r2 6 7 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1490
r3 4 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0980 $X2=0.3510 $Y2=0.1350
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r5 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
.ends

.subckt PM_AO333x2_ASAP7_75t_R%A2 VSS 8 3 4 1
c1 1 VSS 0.0066875f
c2 3 VSS 0.0464558f
c3 4 VSS 0.00500304f
r1 8 7 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1865 $X2=0.2430 $Y2=0.1650
r2 6 7 6.99569 $w=1.3e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1650
r3 4 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0980 $X2=0.2430 $Y2=0.1350
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r5 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AO333x2_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.0424802f
.ends

.subckt PM_AO333x2_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.0423966f
.ends

.subckt PM_AO333x2_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.00475565f
.ends

.subckt PM_AO333x2_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.00461304f
.ends

.subckt PM_AO333x2_ASAP7_75t_R%C3 VSS 8 3 4 1
c1 1 VSS 0.00750045f
c2 3 VSS 0.0465617f
c3 4 VSS 0.00482157f
r1 9 10 6.99569 $w=1.3e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1050 $X2=0.5130 $Y2=0.1350
r2 8 9 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0835 $X2=0.5130 $Y2=0.1050
r3 8 4 1.63233 $w=1.3e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0835 $X2=0.5130 $Y2=0.0765
r4 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r5 1 10 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.1350
+ $X2=0.5130 $Y2=0.1350
.ends

.subckt PM_AO333x2_ASAP7_75t_R%B1 VSS 10 3 4 1
c1 1 VSS 0.00844557f
c2 3 VSS 0.0469442f
c3 4 VSS 0.00525587f
r1 10 9 1.39914 $w=1.3e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1555 $X2=0.4590 $Y2=0.1495
r2 8 9 3.38125 $w=1.3e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1495
r3 4 8 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0980 $X2=0.4590 $Y2=0.1350
r4 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1350
+ $X2=0.4590 $Y2=0.1350
.ends

.subckt PM_AO333x2_ASAP7_75t_R%C1 VSS 8 3 1 4
c1 1 VSS 0.00688802f
c2 3 VSS 0.00848242f
c3 4 VSS 0.00415576f
r1 9 10 7.22888 $w=1.3e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1040 $X2=0.6210 $Y2=0.1350
r2 8 9 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0815 $X2=0.6210 $Y2=0.1040
r3 8 4 1.39914 $w=1.3e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0815 $X2=0.6210 $Y2=0.0755
r4 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1350
r5 1 10 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6210 $Y=0.1350
+ $X2=0.6210 $Y2=0.1350
.ends

.subckt PM_AO333x2_ASAP7_75t_R%C2 VSS 10 3 1 4
c1 1 VSS 0.00630614f
c2 3 VSS 0.00926207f
c3 4 VSS 0.00410343f
r1 10 9 1.16595 $w=1.3e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1535 $X2=0.5670 $Y2=0.1485
r2 8 9 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1485
r3 4 8 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0980 $X2=0.5670 $Y2=0.1350
r4 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1350
+ $X2=0.5670 $Y2=0.1350
.ends

.subckt PM_AO333x2_ASAP7_75t_R%B2 VSS 8 3 4 1
c1 1 VSS 0.00710177f
c2 3 VSS 0.00970554f
c3 4 VSS 0.00473753f
r1 9 10 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1055 $X2=0.4050 $Y2=0.1350
r2 8 9 4.89699 $w=1.3e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0845 $X2=0.4050 $Y2=0.1055
r3 8 4 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0845 $X2=0.4050 $Y2=0.0770
r4 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r5 1 10 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
.ends

.subckt PM_AO333x2_ASAP7_75t_R%Y VSS 24 18 19 33 34 7 2 12 9 10 15 1 8
c1 1 VSS 0.00861726f
c2 2 VSS 0.010614f
c3 7 VSS 0.00455779f
c4 8 VSS 0.00454042f
c5 9 VSS 0.00471211f
c6 10 VSS 0.00241013f
c7 11 VSS 0.0100571f
c8 12 VSS 0.00208451f
c9 13 VSS 0.00137902f
c10 14 VSS 0.00344315f
c11 15 VSS 0.000913771f
r1 34 32 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r2 2 32 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r4 33 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
r5 2 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.2340
r6 28 29 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.0830
+ $Y=0.2340 $X2=0.1080 $Y2=0.2340
r7 11 14 4.06404 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0515 $Y=0.2340 $X2=0.0270 $Y2=0.2340
r8 11 28 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0515
+ $Y=0.2340 $X2=0.0830 $Y2=0.2340
r9 14 27 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0270 $Y2=0.2125
r10 26 27 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1720 $X2=0.0270 $Y2=0.2125
r11 25 26 6.99569 $w=1.3e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1420 $X2=0.0270 $Y2=0.1720
r12 24 25 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1395 $X2=0.0270 $Y2=0.1420
r13 24 23 1.63233 $w=1.3e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1395 $X2=0.0270 $Y2=0.1325
r14 9 13 3.59766 $w=1.692e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1125 $X2=0.0270 $Y2=0.0900
r15 9 23 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1125 $X2=0.0270 $Y2=0.1325
r16 13 22 4.06404 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0900 $X2=0.0515 $Y2=0.0900
r17 10 15 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.0830
+ $Y=0.0900 $X2=0.1080 $Y2=0.0900
r18 10 22 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0830
+ $Y=0.0900 $X2=0.0515 $Y2=0.0900
r19 15 21 1.26576 $w=2.0056e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0900 $X2=0.1080 $Y2=0.0775
r20 20 21 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0650 $X2=0.1080 $Y2=0.0775
r21 12 20 3.38125 $w=1.3e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0505 $X2=0.1080 $Y2=0.0650
r22 1 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1080 $Y2=0.0650
r23 19 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r24 1 17 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r25 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r26 18 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.0935 $Y2=0.0675
.ends

.subckt PM_AO333x2_ASAP7_75t_R%NET22 VSS 16 17 37 38 41 42 13 11 3 12 2 10 1
c1 1 VSS 0.00289997f
c2 2 VSS 0.00318059f
c3 3 VSS 0.00275004f
c4 10 VSS 0.00213512f
c5 11 VSS 0.00210868f
c6 12 VSS 0.0021247f
c7 13 VSS 0.00310906f
r1 42 40 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.2025 $X2=0.6085 $Y2=0.2025
r2 3 40 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.2025 $X2=0.6085 $Y2=0.2025
r3 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2025 $X2=0.5940 $Y2=0.2025
r4 41 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.2025 $X2=0.5795 $Y2=0.2025
r5 38 36 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r6 2 36 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r7 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4860 $Y2=0.2025
r8 37 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r9 3 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2025
+ $X2=0.5940 $Y2=0.1980
r10 2 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2025
+ $X2=0.4860 $Y2=0.1980
r11 31 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5805
+ $Y=0.1980 $X2=0.5940 $Y2=0.1980
r12 30 31 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1980 $X2=0.5805 $Y2=0.1980
r13 29 30 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.5415
+ $Y=0.1980 $X2=0.5670 $Y2=0.1980
r14 28 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5235
+ $Y=0.1980 $X2=0.5415 $Y2=0.1980
r15 27 28 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1980 $X2=0.5235 $Y2=0.1980
r16 26 27 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4995
+ $Y=0.1980 $X2=0.5130 $Y2=0.1980
r17 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.1980 $X2=0.4995 $Y2=0.1980
r18 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4725
+ $Y=0.1980 $X2=0.4860 $Y2=0.1980
r19 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1980 $X2=0.4725 $Y2=0.1980
r20 22 23 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4495
+ $Y=0.1980 $X2=0.4590 $Y2=0.1980
r21 21 22 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4315
+ $Y=0.1980 $X2=0.4495 $Y2=0.1980
r22 20 21 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1980 $X2=0.4315 $Y2=0.1980
r23 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3915
+ $Y=0.1980 $X2=0.4050 $Y2=0.1980
r24 18 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.1980 $X2=0.3915 $Y2=0.1980
r25 13 18 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3665
+ $Y=0.1980 $X2=0.3780 $Y2=0.1980
r26 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.1980
r27 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r28 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r29 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3780 $Y2=0.2025
r30 16 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
.ends

.subckt PM_AO333x2_ASAP7_75t_R%NET40 VSS 16 17 77 78 84 91 94 95 22 1 24 23 28
+ 18 4 5 20 26 6 21 7 19 27 25
c1 1 VSS 0.00818691f
c2 4 VSS 0.00595868f
c3 5 VSS 0.00475714f
c4 6 VSS 0.00599661f
c5 7 VSS 0.00550364f
c6 16 VSS 0.080769f
c7 17 VSS 0.0806685f
c8 18 VSS 0.00434825f
c9 19 VSS 0.00420748f
c10 20 VSS 0.00358783f
c11 21 VSS 0.00384902f
c12 22 VSS 0.00164888f
c13 23 VSS 0.00260996f
c14 24 VSS 0.0483534f
c15 25 VSS 0.0129314f
c16 26 VSS 0.00575935f
c17 27 VSS 0.00257163f
c18 28 VSS 0.000320949f
c19 29 VSS 0.00350091f
c20 30 VSS 0.00316722f
r1 95 93 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r2 5 93 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5400 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r3 20 5 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.2025 $X2=0.5400 $Y2=0.2025
r4 94 20 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.2025 $X2=0.5255 $Y2=0.2025
r5 21 7 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.2025 $X2=0.6460 $Y2=0.2025
r6 91 21 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.2025 $X2=0.6335 $Y2=0.2025
r7 5 88 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.2025
+ $X2=0.5400 $Y2=0.2340
r8 7 85 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.2025
+ $X2=0.6480 $Y2=0.2340
r9 88 89 11.5429 $w=1.3e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.2340 $X2=0.5895 $Y2=0.2340
r10 85 86 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6480
+ $Y=0.2340 $X2=0.6615 $Y2=0.2340
r11 25 85 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6345
+ $Y=0.2340 $X2=0.6480 $Y2=0.2340
r12 25 89 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.6345
+ $Y=0.2340 $X2=0.5895 $Y2=0.2340
r13 30 82 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.2340 $X2=0.6750 $Y2=0.2160
r14 30 86 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6750 $Y=0.2340 $X2=0.6615 $Y2=0.2340
r15 19 6 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0675 $X2=0.6460 $Y2=0.0675
r16 84 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.0675 $X2=0.6335 $Y2=0.0675
r17 81 82 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1980 $X2=0.6750 $Y2=0.2160
r18 80 81 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1765 $X2=0.6750 $Y2=0.1980
r19 79 80 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1170 $X2=0.6750 $Y2=0.1765
r20 26 29 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6750 $Y=0.0575 $X2=0.6750 $Y2=0.0360
r21 26 79 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.0575 $X2=0.6750 $Y2=0.1170
r22 78 76 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r23 4 76 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r24 18 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3240 $Y2=0.0675
r25 77 18 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r26 6 73 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.0675
+ $X2=0.6480 $Y2=0.0360
r27 29 74 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6750 $Y=0.0360 $X2=0.6615 $Y2=0.0360
r28 4 58 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0675
+ $X2=0.3240 $Y2=0.0360
r29 73 74 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6480
+ $Y=0.0360 $X2=0.6615 $Y2=0.0360
r30 72 73 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6345
+ $Y=0.0360 $X2=0.6480 $Y2=0.0360
r31 71 72 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0360 $X2=0.6345 $Y2=0.0360
r32 70 71 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0360 $X2=0.6210 $Y2=0.0360
r33 69 70 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0360 $X2=0.5940 $Y2=0.0360
r34 68 69 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.0360 $X2=0.5670 $Y2=0.0360
r35 67 68 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0360 $X2=0.5400 $Y2=0.0360
r36 66 67 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.0360 $X2=0.5130 $Y2=0.0360
r37 65 66 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0360 $X2=0.4860 $Y2=0.0360
r38 64 65 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4590 $Y2=0.0360
r39 63 64 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r40 62 63 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3800
+ $Y=0.0360 $X2=0.4050 $Y2=0.0360
r41 61 62 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3620
+ $Y=0.0360 $X2=0.3800 $Y2=0.0360
r42 60 61 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0360 $X2=0.3620 $Y2=0.0360
r43 59 60 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.0360 $X2=0.3510 $Y2=0.0360
r44 58 59 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.0360 $X2=0.3375 $Y2=0.0360
r45 57 58 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3105
+ $Y=0.0360 $X2=0.3240 $Y2=0.0360
r46 56 57 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.3105 $Y2=0.0360
r47 55 56 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.2970 $Y2=0.0360
r48 54 55 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r49 53 54 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2180
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r50 52 53 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2000
+ $Y=0.0360 $X2=0.2180 $Y2=0.0360
r51 51 52 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.2000 $Y2=0.0360
r52 24 27 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1710
+ $Y=0.0360 $X2=0.1530 $Y2=0.0360
r53 24 51 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1710
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r54 27 50 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1530 $Y=0.0360 $X2=0.1530 $Y2=0.0575
r55 49 50 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1530
+ $Y=0.0845 $X2=0.1530 $Y2=0.0575
r56 23 28 3.59766 $w=1.692e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1530 $Y=0.1125 $X2=0.1530 $Y2=0.1350
r57 23 49 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1530
+ $Y=0.1125 $X2=0.1530 $Y2=0.0845
r58 28 47 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1530
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r59 17 40 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1350 $Y2=0.1350
r60 46 47 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1240
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r61 45 46 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1195
+ $Y=0.1350 $X2=0.1240 $Y2=0.1350
r62 44 45 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.1035
+ $Y=0.1350 $X2=0.1195 $Y2=0.1350
r63 43 44 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.1035 $Y2=0.1350
r64 22 43 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0695
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r65 40 47 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
r66 39 40 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1255
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r67 37 39 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1350 $X2=0.1255 $Y2=0.1350
r68 36 37 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1350 $X2=0.1225 $Y2=0.1350
r69 35 36 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1350 $X2=0.1080 $Y2=0.1350
r70 33 35 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0905 $Y=0.1350 $X2=0.0935 $Y2=0.1350
r71 32 33 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0905 $Y2=0.1350
r72 32 43 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
r73 1 32 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r74 1 34 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1350 $X2=0.0705 $Y2=0.1350
r75 16 32 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0810 $Y2=0.1350
r76 16 34 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.0810 $Y=0.1350 $X2=0.0705 $Y2=0.1350
r77 16 35 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1350
.ends


*
.SUBCKT AO333x2_ASAP7_75t_R VSS VDD A3 A2 A1 B3 B2 B1 C3 C2 C1 Y
*
* VSS VSS
* VDD VDD
* A3 A3
* A2 A2
* A1 A1
* B3 B3
* B2 B2
* B1 B1
* C3 C3
* C2 C2
* C1 C1
* Y Y
*
*

MM3 N_MM3_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3@2 N_MM3@2_d N_MM4@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM19 N_MM19_d N_MM17_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM18 N_MM18_d N_MM16_g N_MM18_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM14 N_MM14_d N_MM15_g N_MM14_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM13_g N_MM10_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM12_g N_MM9_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM5_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM6_g N_MM1_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM0_g N_MM0_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@2 N_MM4@2_d N_MM4@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM17 N_MM17_d N_MM17_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM16 N_MM16_d N_MM16_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM15 N_MM15_d N_MM15_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM13 N_MM13_d N_MM13_g N_MM13_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM12 N_MM12_d N_MM12_g N_MM12_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 N_MM11_d N_MM11_g N_MM11_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM6_g N_MM6_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM0_g N_MM7_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AO333x2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AO333x2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AO333x2_ASAP7_75t_R%NET54 VSS N_MM2_d N_MM1_s N_NET54_1
+ PM_AO333x2_ASAP7_75t_R%NET54
cc_1 N_NET54_1 N_MM5_g 0.0173884f
cc_2 N_NET54_1 N_MM6_g 0.0173089f
x_PM_AO333x2_ASAP7_75t_R%NET55 VSS N_MM0_s N_MM1_d N_NET55_1
+ PM_AO333x2_ASAP7_75t_R%NET55
cc_3 N_NET55_1 N_MM6_g 0.0174376f
cc_4 N_NET55_1 N_MM0_g 0.0172824f
x_PM_AO333x2_ASAP7_75t_R%NET59 VSS N_MM18_d N_MM14_s N_NET59_1
+ PM_AO333x2_ASAP7_75t_R%NET59
cc_5 N_NET59_1 N_MM16_g 0.0174209f
cc_6 N_NET59_1 N_MM15_g 0.0172753f
x_PM_AO333x2_ASAP7_75t_R%NET57 VSS N_MM9_s N_MM8_d N_NET57_1
+ PM_AO333x2_ASAP7_75t_R%NET57
cc_7 N_NET57_1 N_MM12_g 0.0174078f
cc_8 N_NET57_1 N_MM11_g 0.0173048f
x_PM_AO333x2_ASAP7_75t_R%NET56 VSS N_MM10_s N_MM9_d N_NET56_1
+ PM_AO333x2_ASAP7_75t_R%NET56
cc_9 N_NET56_1 N_MM13_g 0.0173598f
cc_10 N_NET56_1 N_MM12_g 0.0173217f
x_PM_AO333x2_ASAP7_75t_R%NET58 VSS N_MM19_d N_MM18_s N_NET58_1
+ PM_AO333x2_ASAP7_75t_R%NET58
cc_11 N_NET58_1 N_MM17_g 0.0173435f
cc_12 N_NET58_1 N_MM16_g 0.0173545f
x_PM_AO333x2_ASAP7_75t_R%NET24 VSS N_MM17_d N_MM16_d N_MM15_d N_MM13_s N_MM12_s
+ N_MM11_s N_NET24_1 N_NET24_10 N_NET24_13 N_NET24_2 N_NET24_11 N_NET24_12
+ N_NET24_3 PM_AO333x2_ASAP7_75t_R%NET24
cc_13 N_NET24_1 N_A3_4 0.00106067f
cc_14 N_NET24_1 N_MM17_g 0.00117681f
cc_15 N_NET24_10 N_MM17_g 0.034716f
cc_16 N_NET24_10 N_A2_1 0.00066572f
cc_17 N_NET24_13 N_A2_4 0.00108082f
cc_18 N_NET24_1 N_MM16_g 0.00117006f
cc_19 N_NET24_1 N_A2_4 0.00162162f
cc_20 N_NET24_10 N_MM16_g 0.0334311f
cc_21 N_NET24_13 N_A1_4 0.00115938f
cc_22 N_NET24_2 N_MM15_g 0.0011692f
cc_23 N_NET24_2 N_A1_4 0.00168803f
cc_24 N_NET24_11 N_MM15_g 0.0342236f
cc_25 N_NET24_11 N_B3_1 0.000724565f
cc_26 N_NET24_2 N_MM13_g 0.000918653f
cc_27 N_NET24_11 N_MM13_g 0.0338718f
cc_28 N_NET24_12 N_B2_1 0.00065993f
cc_29 N_NET24_3 N_MM12_g 0.0009101f
cc_30 N_NET24_12 N_MM12_g 0.0336627f
cc_31 N_NET24_12 N_B1_1 0.000674321f
cc_32 N_NET24_3 N_MM11_g 0.000899941f
cc_33 N_NET24_12 N_MM11_g 0.0334195f
x_PM_AO333x2_ASAP7_75t_R%A3 VSS A3 N_MM17_g N_A3_4 N_A3_1
+ PM_AO333x2_ASAP7_75t_R%A3
cc_34 N_A3_4 N_NET40_22 0.000305096f
cc_35 N_A3_4 N_NET40_1 0.000305646f
cc_36 N_A3_1 N_NET40_1 0.000978751f
cc_37 N_A3_4 N_NET40_24 0.00104055f
cc_38 N_A3_4 N_NET40_23 0.00221644f
cc_39 N_MM17_g N_MM4@2_g 0.00339746f
cc_40 N_A3_4 N_NET40_28 0.0064746f
x_PM_AO333x2_ASAP7_75t_R%A1 VSS A1 N_MM15_g N_A1_1 N_A1_4
+ PM_AO333x2_ASAP7_75t_R%A1
cc_41 N_MM15_g N_NET40_4 0.00180486f
cc_42 N_A1_1 N_NET40_18 0.000880955f
cc_43 N_A1_4 N_NET40_24 0.00133784f
cc_44 N_A1_4 N_NET40_4 0.00186408f
cc_45 N_MM15_g N_NET40_18 0.0355407f
cc_46 N_A1_1 N_A2_1 0.0013377f
cc_47 N_A1_4 N_A2_4 0.00476599f
cc_48 N_MM15_g N_MM16_g 0.00615893f
x_PM_AO333x2_ASAP7_75t_R%B3 VSS B3 N_MM13_g N_B3_1 N_B3_4
+ PM_AO333x2_ASAP7_75t_R%B3
cc_49 N_MM13_g N_NET40_4 0.00179374f
cc_50 N_B3_1 N_NET40_18 0.000919135f
cc_51 N_B3_4 N_NET40_24 0.00130191f
cc_52 N_B3_4 N_NET40_4 0.00176322f
cc_53 N_MM13_g N_NET40_18 0.0354088f
cc_54 N_B3_1 N_A1_4 0.000941972f
cc_55 N_MM13_g N_MM15_g 0.00327896f
cc_56 N_B3_4 N_A1_4 0.00437288f
x_PM_AO333x2_ASAP7_75t_R%A2 VSS A2 N_MM16_g N_A2_4 N_A2_1
+ PM_AO333x2_ASAP7_75t_R%A2
cc_57 N_A2_4 N_NET40_23 8.39341e-20
cc_58 N_A2_4 N_NET40_18 0.000666603f
cc_59 N_A2_4 N_NET40_4 0.000275677f
cc_60 N_A2_4 N_NET40_24 0.00143466f
cc_61 N_A2_4 N_NET40_28 0.00184955f
cc_62 N_A2_1 N_A3_1 0.00137236f
cc_63 N_A2_4 N_A3_4 0.0049341f
cc_64 N_MM16_g N_MM17_g 0.00621702f
x_PM_AO333x2_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_AO333x2_ASAP7_75t_R%noxref_22
cc_65 N_noxref_22_1 N_MM3_g 0.00149695f
cc_66 N_noxref_22_1 N_Y_7 0.000700363f
x_PM_AO333x2_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_AO333x2_ASAP7_75t_R%noxref_23
cc_67 N_noxref_23_1 N_MM3_g 0.00149326f
cc_68 N_noxref_23_1 N_Y_8 0.00081649f
cc_69 N_noxref_23_1 N_noxref_22_1 0.00177611f
x_PM_AO333x2_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_AO333x2_ASAP7_75t_R%noxref_24
cc_70 N_noxref_24_1 N_NET40_21 8.86546e-20
cc_71 N_noxref_24_1 N_NET40_26 0.000322451f
cc_72 N_noxref_24_1 N_NET40_6 0.000506288f
cc_73 N_noxref_24_1 N_NET40_19 0.0375451f
cc_74 N_noxref_24_1 N_MM0_g 0.00146219f
x_PM_AO333x2_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_AO333x2_ASAP7_75t_R%noxref_25
cc_75 N_noxref_25_1 N_NET40_19 8.95035e-20
cc_76 N_noxref_25_1 N_NET40_26 0.000321983f
cc_77 N_noxref_25_1 N_NET40_7 0.000503616f
cc_78 N_noxref_25_1 N_NET40_21 0.0376255f
cc_79 N_noxref_25_1 N_MM0_g 0.00144534f
cc_80 N_noxref_25_1 N_noxref_24_1 0.0017751f
x_PM_AO333x2_ASAP7_75t_R%C3 VSS C3 N_MM5_g N_C3_4 N_C3_1
+ PM_AO333x2_ASAP7_75t_R%C3
cc_81 N_MM5_g N_NET40_5 0.00115836f
cc_82 N_C3_4 N_NET40_24 0.0013707f
cc_83 N_C3_4 N_NET40_5 0.00152587f
cc_84 N_MM5_g N_NET40_20 0.0355202f
cc_85 N_C3_1 N_B1_1 0.000971352f
cc_86 N_C3_4 N_B1_4 0.00321659f
cc_87 N_MM5_g N_MM11_g 0.00402371f
x_PM_AO333x2_ASAP7_75t_R%B1 VSS B1 N_MM11_g N_B1_4 N_B1_1
+ PM_AO333x2_ASAP7_75t_R%B1
cc_88 N_B1_4 N_NET40_24 0.00303412f
cc_89 N_B1_1 N_B2_1 0.00138709f
cc_90 N_B1_4 N_B2_4 0.00333516f
cc_91 N_MM11_g N_MM12_g 0.00608167f
x_PM_AO333x2_ASAP7_75t_R%C1 VSS C1 N_MM0_g N_C1_1 N_C1_4
+ PM_AO333x2_ASAP7_75t_R%C1
cc_92 N_MM0_g N_NET40_6 0.00186403f
cc_93 N_MM0_g N_NET40_21 0.0158857f
cc_94 N_C1_1 N_NET40_7 0.000783432f
cc_95 N_MM0_g N_NET40_7 0.00107661f
cc_96 N_C1_4 N_NET40_24 0.00123191f
cc_97 N_C1_1 N_NET40_21 0.00171839f
cc_98 N_C1_4 N_NET40_26 0.00605515f
cc_99 N_MM0_g N_NET40_19 0.0547221f
cc_100 N_C1_1 N_C2_1 0.00125572f
cc_101 N_C1_4 N_C2_4 0.00336323f
cc_102 N_MM0_g N_MM6_g 0.00597343f
x_PM_AO333x2_ASAP7_75t_R%C2 VSS C2 N_MM6_g N_C2_1 N_C2_4
+ PM_AO333x2_ASAP7_75t_R%C2
cc_103 N_MM6_g N_NET40_26 0.000130921f
cc_104 N_MM6_g N_NET40_6 0.000272382f
cc_105 N_MM6_g N_NET40_5 0.00124485f
cc_106 N_C2_1 N_NET40_20 0.000827813f
cc_107 N_C2_4 N_NET40_24 0.00144997f
cc_108 N_C2_4 N_NET40_5 0.00167007f
cc_109 N_MM6_g N_NET40_20 0.0352614f
cc_110 N_C2_1 N_C3_1 0.00133047f
cc_111 N_C2_4 N_C3_4 0.0034115f
cc_112 N_MM6_g N_MM5_g 0.00605593f
x_PM_AO333x2_ASAP7_75t_R%B2 VSS B2 N_MM12_g N_B2_4 N_B2_1
+ PM_AO333x2_ASAP7_75t_R%B2
cc_113 N_B2_4 N_NET40_18 0.000541359f
cc_114 N_B2_4 N_NET40_4 0.000277803f
cc_115 N_B2_4 N_NET40_24 0.00316178f
cc_116 N_B2_1 N_B3_1 0.00144986f
cc_117 N_B2_4 N_B3_4 0.0036171f
cc_118 N_MM12_g N_MM13_g 0.00596385f
x_PM_AO333x2_ASAP7_75t_R%Y VSS Y N_MM3_d N_MM3@2_d N_MM4_d N_MM4@2_d N_Y_7
+ N_Y_2 N_Y_12 N_Y_9 N_Y_10 N_Y_15 N_Y_1 N_Y_8 PM_AO333x2_ASAP7_75t_R%Y
cc_119 N_Y_7 N_NET40_28 0.000200589f
cc_120 N_Y_7 N_NET40_23 0.000322758f
cc_121 N_Y_7 N_NET40_27 0.000368986f
cc_122 N_Y_7 N_NET40_22 0.000415154f
cc_123 N_Y_7 N_NET40_1 0.000512025f
cc_124 N_Y_2 N_NET40_1 0.000950244f
cc_125 N_Y_12 N_NET40_23 0.00104875f
cc_126 N_Y_9 N_NET40_22 0.00125033f
cc_127 N_Y_10 N_NET40_22 0.00130788f
cc_128 N_Y_15 N_NET40_23 0.00178806f
cc_129 N_Y_2 N_MM3_g 0.00210612f
cc_130 N_Y_1 N_MM3_g 0.00213977f
cc_131 N_Y_15 N_NET40_22 0.0040065f
cc_132 N_Y_8 N_NET40_1 0.00439206f
cc_133 N_Y_8 N_MM3_g 0.029791f
cc_134 N_Y_7 N_MM4@2_g 0.0369922f
cc_135 N_Y_7 N_MM3_g 0.0688821f
x_PM_AO333x2_ASAP7_75t_R%NET22 VSS N_MM13_d N_MM12_d N_MM11_d N_MM5_s N_MM6_s
+ N_MM7_s N_NET22_13 N_NET22_11 N_NET22_3 N_NET22_12 N_NET22_2 N_NET22_10
+ N_NET22_1 PM_AO333x2_ASAP7_75t_R%NET22
cc_136 N_NET22_13 N_NET40_20 9.70111e-20
cc_137 N_NET22_13 N_NET40_5 0.00094042f
cc_138 N_NET22_13 N_NET40_7 0.000300289f
cc_139 N_NET22_13 N_NET40_21 0.000555378f
cc_140 N_NET22_11 N_NET40_20 0.00167036f
cc_141 N_NET22_13 N_NET40_26 0.000632744f
cc_142 N_NET22_3 N_NET40_25 0.000656501f
cc_143 N_NET22_12 N_NET40_20 0.00111355f
cc_144 N_NET22_3 N_NET40_7 0.00144399f
cc_145 N_NET22_3 N_NET40_5 0.00278014f
cc_146 N_NET22_2 N_NET40_5 0.00427708f
cc_147 N_NET22_13 N_NET40_25 0.0106047f
cc_148 N_NET22_10 N_B3_1 0.000726745f
cc_149 N_NET22_1 N_B3_4 0.00076553f
cc_150 N_NET22_1 N_MM13_g 0.000848325f
cc_151 N_NET22_10 N_MM13_g 0.0340503f
cc_152 N_NET22_10 N_B2_1 0.00073835f
cc_153 N_NET22_1 N_MM12_g 0.00087943f
cc_154 N_NET22_13 N_B2_4 0.00119463f
cc_155 N_NET22_1 N_B2_4 0.00123945f
cc_156 N_NET22_10 N_MM12_g 0.0335058f
cc_157 N_NET22_11 N_B1_1 0.000683946f
cc_158 N_NET22_2 N_MM11_g 0.000877827f
cc_159 N_NET22_13 N_B1_4 0.00121857f
cc_160 N_NET22_2 N_B1_4 0.00123591f
cc_161 N_NET22_11 N_MM11_g 0.0335773f
cc_162 N_NET22_2 N_MM5_g 0.000876702f
cc_163 N_NET22_13 N_C3_4 0.00121065f
cc_164 N_NET22_2 N_C3_4 0.00125597f
cc_165 N_NET22_11 N_MM5_g 0.0341756f
cc_166 N_NET22_12 N_C2_1 0.00069779f
cc_167 N_NET22_3 N_MM6_g 0.000871049f
cc_168 N_NET22_3 N_C2_4 0.00121262f
cc_169 N_NET22_13 N_C2_4 0.00123982f
cc_170 N_NET22_12 N_MM6_g 0.0336353f
cc_171 N_NET22_12 N_C1_1 0.0006938f
cc_172 N_NET22_3 N_MM0_g 0.000892694f
cc_173 N_NET22_13 N_C1_4 0.000907661f
cc_174 N_NET22_3 N_C1_4 0.000962843f
cc_175 N_NET22_12 N_MM0_g 0.0334821f
cc_176 N_NET22_10 N_NET24_13 0.000554959f
cc_177 N_NET22_13 N_NET24_3 0.000651194f
cc_178 N_NET22_1 N_NET24_13 0.000705163f
cc_179 N_NET22_10 N_NET24_11 0.00111658f
cc_180 N_NET22_10 N_NET24_12 0.00111986f
cc_181 N_NET22_2 N_NET24_3 0.00124193f
cc_182 N_NET22_1 N_NET24_3 0.00301376f
cc_183 N_NET22_1 N_NET24_2 0.00410421f
cc_184 N_NET22_13 N_NET24_13 0.0100848f
x_PM_AO333x2_ASAP7_75t_R%NET40 VSS N_MM3_g N_MM4@2_g N_MM14_d N_MM10_d N_MM0_d
+ N_MM7_d N_MM5_d N_MM6_d N_NET40_22 N_NET40_1 N_NET40_24 N_NET40_23 N_NET40_28
+ N_NET40_18 N_NET40_4 N_NET40_5 N_NET40_20 N_NET40_26 N_NET40_6 N_NET40_21
+ N_NET40_7 N_NET40_19 N_NET40_27 N_NET40_25 PM_AO333x2_ASAP7_75t_R%NET40
*END of AO333x2_ASAP7_75t_R.pxi
.ENDS
** Design:	AO33x2_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AO33x2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AO33x2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AO33x2_ASAP7_75t_R%NET40 VSS 2 3 1
c1 1 VSS 0.000964898f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2700 $Y2=0.0675
.ends

.subckt PM_AO33x2_ASAP7_75t_R%NET024 VSS 2 3 1
c1 1 VSS 0.000934274f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2160 $Y2=0.0675
.ends

.subckt PM_AO33x2_ASAP7_75t_R%NET39 VSS 2 3 1
c1 1 VSS 0.000954705f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3780 $Y2=0.0675
.ends

.subckt PM_AO33x2_ASAP7_75t_R%NET022 VSS 2 3 1
c1 1 VSS 0.000939443f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4320 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4320 $Y2=0.0675
.ends

.subckt PM_AO33x2_ASAP7_75t_R%A1 VSS 6 3 1 4
c1 1 VSS 0.0065239f
c2 3 VSS 0.0418016f
c3 4 VSS 0.00464566f
r1 7 8 3.20636 $w=1.3e-08 $l=1.38e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1212 $X2=0.2970 $Y2=0.1350
r2 6 7 1.22425 $w=1.3e-08 $l=5.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1160 $X2=0.2970 $Y2=0.1212
r3 6 4 5.42166 $w=1.3e-08 $l=2.33e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1160 $X2=0.2970 $Y2=0.0927
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_AO33x2_ASAP7_75t_R%A2 VSS 8 3 4 1
c1 1 VSS 0.00563028f
c2 3 VSS 0.0423632f
c3 4 VSS 0.00423411f
r1 8 7 5.42166 $w=1.3e-08 $l=2.33e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1900 $X2=0.2430 $Y2=0.1667
r2 6 7 7.40378 $w=1.3e-08 $l=3.17e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1667
r3 4 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0980 $X2=0.2430 $Y2=0.1350
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r5 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AO33x2_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.042388f
.ends

.subckt PM_AO33x2_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.00483087f
.ends

.subckt PM_AO33x2_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.0419736f
.ends

.subckt PM_AO33x2_ASAP7_75t_R%A3 VSS 8 3 4 1
c1 1 VSS 0.00711405f
c2 3 VSS 0.083482f
c3 4 VSS 0.00621274f
r1 8 7 0.349785 $w=1.3e-08 $l=1.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1465 $X2=0.1890 $Y2=0.1450
r2 6 7 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1450
r3 4 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0980 $X2=0.1890 $Y2=0.1350
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r5 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AO33x2_ASAP7_75t_R%Y VSS 25 17 18 33 34 7 8 9 2 1 14
c1 1 VSS 0.00904408f
c2 2 VSS 0.0105543f
c3 7 VSS 0.00458638f
c4 8 VSS 0.00455981f
c5 9 VSS 0.0053691f
c6 10 VSS 0.00277094f
c7 11 VSS 0.00954301f
c8 12 VSS 0.00153546f
c9 13 VSS 0.00338781f
c10 14 VSS 0.0033827f
r1 34 32 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r2 2 32 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r4 33 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
r5 2 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.2340
r6 28 29 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.0830
+ $Y=0.2340 $X2=0.1080 $Y2=0.2340
r7 11 13 4.06404 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0515 $Y=0.2340 $X2=0.0270 $Y2=0.2340
r8 11 28 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0515
+ $Y=0.2340 $X2=0.0830 $Y2=0.2340
r9 13 27 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0270 $Y2=0.2125
r10 26 27 9.0944 $w=1.3e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1735 $X2=0.0270 $Y2=0.2125
r11 25 26 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1465 $X2=0.0270 $Y2=0.1735
r12 25 24 0.349785 $w=1.3e-08 $l=1.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1465 $X2=0.0270 $Y2=0.1450
r13 23 24 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1350 $X2=0.0270 $Y2=0.1450
r14 9 12 5.11339 $w=1.60414e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1060 $X2=0.0270 $Y2=0.0770
r15 9 23 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1060 $X2=0.0270 $Y2=0.1350
r16 12 22 4.06404 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0770 $X2=0.0515 $Y2=0.0770
r17 10 21 4.64944 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.0830
+ $Y=0.0770 $X2=0.1080 $Y2=0.0770
r18 10 22 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0830
+ $Y=0.0770 $X2=0.0515 $Y2=0.0770
r19 20 21 1.50137 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0655 $X2=0.1080 $Y2=0.0770
r20 19 20 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0540 $X2=0.1080 $Y2=0.0655
r21 14 19 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0410 $X2=0.1080 $Y2=0.0540
r22 1 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1080 $Y2=0.0540
r23 18 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r24 1 16 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r25 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r26 17 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.0935 $Y2=0.0675
.ends

.subckt PM_AO33x2_ASAP7_75t_R%B1 VSS 6 3 1 4
c1 1 VSS 0.00546724f
c2 3 VSS 0.00800036f
c3 4 VSS 0.00367847f
r1 7 8 7.46207 $w=1.3e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1030 $X2=0.3510 $Y2=0.1350
r2 6 7 5.47996 $w=1.3e-08 $l=2.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0795 $X2=0.3510 $Y2=0.1030
r3 6 4 1.16595 $w=1.3e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0795 $X2=0.3510 $Y2=0.0745
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
.ends

.subckt PM_AO33x2_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.0423805f
.ends

.subckt PM_AO33x2_ASAP7_75t_R%B3 VSS 8 3 1 4
c1 1 VSS 0.00621305f
c2 3 VSS 0.0458647f
c3 4 VSS 0.00401628f
r1 8 7 0.349785 $w=1.3e-08 $l=1.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1465 $X2=0.4590 $Y2=0.1450
r2 6 7 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1450
r3 4 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0980 $X2=0.4590 $Y2=0.1350
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r5 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1350
+ $X2=0.4590 $Y2=0.1350
.ends

.subckt PM_AO33x2_ASAP7_75t_R%B2 VSS 8 3 1 4
c1 1 VSS 0.00490002f
c2 3 VSS 0.00861951f
c3 4 VSS 0.00345013f
r1 8 7 0.349785 $w=1.3e-08 $l=1.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1465 $X2=0.4050 $Y2=0.1450
r2 6 7 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1450
r3 4 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0980 $X2=0.4050 $Y2=0.1350
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r5 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
.ends

.subckt PM_AO33x2_ASAP7_75t_R%NET15 VSS 16 17 33 34 37 38 13 11 3 12 2 1 10
c1 1 VSS 0.0102509f
c2 2 VSS 0.00701053f
c3 3 VSS 0.00457429f
c4 10 VSS 0.00449966f
c5 11 VSS 0.00321213f
c6 12 VSS 0.00210444f
c7 13 VSS 0.0212992f
r1 38 36 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2160 $X2=0.4465 $Y2=0.2160
r2 3 36 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2160 $X2=0.4465 $Y2=0.2160
r3 12 3 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2160 $X2=0.4320 $Y2=0.2160
r4 37 12 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2160 $X2=0.4175 $Y2=0.2160
r5 34 32 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2160 $X2=0.3385 $Y2=0.2160
r6 2 32 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2160 $X2=0.3385 $Y2=0.2160
r7 11 2 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2160 $X2=0.3240 $Y2=0.2160
r8 33 11 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2160 $X2=0.3095 $Y2=0.2160
r9 3 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.2340
r10 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.2340
r11 28 29 9.32759 $w=1.3e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3920
+ $Y=0.2340 $X2=0.4320 $Y2=0.2340
r12 27 28 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3605
+ $Y=0.2340 $X2=0.3920 $Y2=0.2340
r13 26 27 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.2340 $X2=0.3605 $Y2=0.2340
r14 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.2340 $X2=0.3510 $Y2=0.2340
r15 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.2340 $X2=0.3375 $Y2=0.2340
r16 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3105
+ $Y=0.2340 $X2=0.3240 $Y2=0.2340
r17 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.2340 $X2=0.3105 $Y2=0.2340
r18 21 22 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.2970 $Y2=0.2340
r19 20 21 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r20 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.2340 $X2=0.2430 $Y2=0.2340
r21 18 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2295 $Y2=0.2340
r22 13 18 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.2030
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r23 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.2340
r24 17 15 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2160 $X2=0.2305 $Y2=0.2160
r25 1 15 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2160 $X2=0.2305 $Y2=0.2160
r26 10 1 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2160 $X2=0.2160 $Y2=0.2160
r27 16 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2160 $X2=0.2015 $Y2=0.2160
.ends

.subckt PM_AO33x2_ASAP7_75t_R%NET020 VSS 12 13 63 64 77 80 81 1 19 18 23 14 3
+ 20 15 4 5 16 21 17 22
c1 1 VSS 0.00764737f
c2 3 VSS 0.00574609f
c3 4 VSS 0.00296285f
c4 5 VSS 0.00482854f
c5 12 VSS 0.0808383f
c6 13 VSS 0.0804378f
c7 14 VSS 0.00482095f
c8 15 VSS 0.00368212f
c9 16 VSS 0.00421227f
c10 17 VSS 0.00197952f
c11 18 VSS 0.00266209f
c12 19 VSS 0.0335102f
c13 20 VSS 0.00300658f
c14 21 VSS 0.00773192f
c15 22 VSS 0.00241216f
c16 23 VSS 0.000340198f
c17 24 VSS 0.00407845f
c18 25 VSS 0.00191952f
r1 81 79 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2160 $X2=0.3925 $Y2=0.2160
r2 4 79 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.2160 $X2=0.3925 $Y2=0.2160
r3 15 4 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2160 $X2=0.3780 $Y2=0.2160
r4 80 15 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2160 $X2=0.3635 $Y2=0.2160
r5 16 5 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2160 $X2=0.4840 $Y2=0.2160
r6 77 16 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2160 $X2=0.4715 $Y2=0.2160
r7 4 74 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.1980
r8 5 67 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2025
+ $X2=0.4860 $Y2=0.1980
r9 74 75 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.1980 $X2=0.3915 $Y2=0.1980
r10 72 75 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1980 $X2=0.3915 $Y2=0.1980
r11 71 72 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.4315
+ $Y=0.1980 $X2=0.4050 $Y2=0.1980
r12 70 71 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4495
+ $Y=0.1980 $X2=0.4315 $Y2=0.1980
r13 69 70 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1980 $X2=0.4495 $Y2=0.1980
r14 67 68 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.1980 $X2=0.4995 $Y2=0.1980
r15 20 67 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4725
+ $Y=0.1980 $X2=0.4860 $Y2=0.1980
r16 20 69 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4725
+ $Y=0.1980 $X2=0.4590 $Y2=0.1980
r17 25 66 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1980 $X2=0.5130 $Y2=0.1765
r18 25 68 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1980 $X2=0.4995 $Y2=0.1980
r19 65 66 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1170 $X2=0.5130 $Y2=0.1765
r20 21 24 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.0575 $X2=0.5130 $Y2=0.0360
r21 21 65 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0575 $X2=0.5130 $Y2=0.1170
r22 64 62 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r23 3 62 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r24 14 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3240 $Y2=0.0675
r25 63 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r26 24 60 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.0360 $X2=0.4860 $Y2=0.0360
r27 3 52 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0675
+ $X2=0.3240 $Y2=0.0360
r28 59 60 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0360 $X2=0.4860 $Y2=0.0360
r29 58 59 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4590 $Y2=0.0360
r30 57 58 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r31 56 57 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.3785
+ $Y=0.0360 $X2=0.4050 $Y2=0.0360
r32 55 56 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3605
+ $Y=0.0360 $X2=0.3785 $Y2=0.0360
r33 54 55 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0360 $X2=0.3605 $Y2=0.0360
r34 53 54 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.0360 $X2=0.3510 $Y2=0.0360
r35 52 53 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.0360 $X2=0.3375 $Y2=0.0360
r36 51 52 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3105
+ $Y=0.0360 $X2=0.3240 $Y2=0.0360
r37 50 51 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.3105 $Y2=0.0360
r38 49 50 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.2970 $Y2=0.0360
r39 48 49 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r40 47 48 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.2165
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r41 46 47 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1985
+ $Y=0.0360 $X2=0.2165 $Y2=0.0360
r42 45 46 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.1985 $Y2=0.0360
r43 19 22 2.50689 $w=1.45385e-08 $l=1.86815e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1710 $Y=0.0360 $X2=0.1530 $Y2=0.0410
r44 19 45 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1710
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r45 22 43 3.32305 $w=1.42121e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1530 $Y=0.0410 $X2=0.1530 $Y2=0.0575
r46 42 43 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1530
+ $Y=0.0780 $X2=0.1530 $Y2=0.0575
r47 18 23 5.11339 $w=1.60414e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1530 $Y=0.1060 $X2=0.1530 $Y2=0.1350
r48 18 42 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1530
+ $Y=0.1060 $X2=0.1530 $Y2=0.0780
r49 23 40 3.01468 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1530
+ $Y=0.1350 $X2=0.1330 $Y2=0.1350
r50 13 34 2.68099 $w=1.25e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1345
r51 39 40 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1195
+ $Y=0.1350 $X2=0.1330 $Y2=0.1350
r52 38 39 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.1350 $X2=0.1195 $Y2=0.1350
r53 37 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.1350 $X2=0.1080 $Y2=0.1350
r54 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0945 $Y2=0.1350
r55 17 36 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0695
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r56 32 34 3.5124 $w=2.166e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1345 $X2=0.1350 $Y2=0.1345
r57 31 32 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1345 $X2=0.1225 $Y2=0.1345
r58 30 31 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1345 $X2=0.1080 $Y2=0.1345
r59 28 30 1.26439 $w=1.74167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0905 $Y=0.1345 $X2=0.0935 $Y2=0.1345
r60 27 28 2.24801 $w=2.3e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0810
+ $Y=0.1345 $X2=0.0905 $Y2=0.1345
r61 27 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1345
+ $X2=0.0810 $Y2=0.1350
r62 1 27 2.24801 $w=2.3e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1345 $X2=0.0810 $Y2=0.1345
r63 1 29 0.347531 $w=1.965e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1345 $X2=0.0705 $Y2=0.1345
r64 12 27 2.44436 $w=1.30368e-07 $l=5e-10 $layer=LIG $thickness=5.22105e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0810 $Y2=0.1345
r65 12 29 0.54388 $w=2.16967e-07 $l=1.05119e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.0810 $Y=0.1350 $X2=0.0705 $Y2=0.1345
r66 12 30 1.46074 $w=1.8486e-07 $l=1.251e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1345
.ends


*
.SUBCKT AO33x2_ASAP7_75t_R VSS VDD A3 A2 A1 B1 B2 B3 Y
*
* VSS VSS
* VDD VDD
* A3 A3
* A2 A2
* A1 A1
* B1 B1
* B2 B2
* B3 B3
* Y Y
*
*

MM24 N_MM24_d N_MM24_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24@2 N_MM24@2_d N_MM24@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM5_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM4_g N_MM0_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM21_g N_MM7_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM2_g N_MM10_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM3_g N_MM8_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM6_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25 N_MM25_d N_MM24_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25@2 N_MM25@2_d N_MM24@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM4 N_MM4_d N_MM4_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM21 N_MM21_d N_MM21_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2 N_MM2_d N_MM2_g N_MM2_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g N_MM3_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM6 N_MM6_d N_MM6_g N_MM6_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2


*include "AO33x2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AO33x2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AO33x2_ASAP7_75t_R%NET40 VSS N_MM0_d N_MM7_s N_NET40_1
+ PM_AO33x2_ASAP7_75t_R%NET40
cc_1 N_NET40_1 N_MM4_g 0.0173445f
cc_2 N_NET40_1 N_MM21_g 0.0174252f
x_PM_AO33x2_ASAP7_75t_R%NET024 VSS N_MM1_d N_MM0_s N_NET024_1
+ PM_AO33x2_ASAP7_75t_R%NET024
cc_3 N_NET024_1 N_MM5_g 0.0173373f
cc_4 N_NET024_1 N_MM4_g 0.0174417f
x_PM_AO33x2_ASAP7_75t_R%NET39 VSS N_MM10_s N_MM8_d N_NET39_1
+ PM_AO33x2_ASAP7_75t_R%NET39
cc_5 N_NET39_1 N_MM2_g 0.0173234f
cc_6 N_NET39_1 N_MM3_g 0.0174555f
x_PM_AO33x2_ASAP7_75t_R%NET022 VSS N_MM8_s N_MM9_d N_NET022_1
+ PM_AO33x2_ASAP7_75t_R%NET022
cc_7 N_NET022_1 N_MM3_g 0.0172287f
cc_8 N_NET022_1 N_MM6_g 0.0172277f
x_PM_AO33x2_ASAP7_75t_R%A1 VSS A1 N_MM21_g N_A1_1 N_A1_4
+ PM_AO33x2_ASAP7_75t_R%A1
cc_9 N_MM21_g N_NET020_20 0.000205667f
cc_10 N_MM21_g N_NET020_3 0.0018039f
cc_11 N_A1_1 N_NET020_14 0.000780932f
cc_12 N_A1_4 N_NET020_19 0.00131034f
cc_13 N_A1_4 N_NET020_3 0.00215178f
cc_14 N_MM21_g N_NET020_14 0.0357682f
cc_15 N_A1_1 N_A2_1 0.00131165f
cc_16 N_A1_4 N_A2_4 0.00484411f
cc_17 N_MM21_g N_MM4_g 0.00727003f
x_PM_AO33x2_ASAP7_75t_R%A2 VSS A2 N_MM4_g N_A2_4 N_A2_1 PM_AO33x2_ASAP7_75t_R%A2
cc_18 N_A2_4 N_NET020_14 0.000121591f
cc_19 N_A2_4 N_NET020_3 0.000276738f
cc_20 N_MM4_g N_NET020_14 0.000447036f
cc_21 N_A2_4 N_NET020_19 0.00141716f
cc_22 N_A2_4 N_NET020_23 0.00197194f
cc_23 N_A2_1 N_A3_1 0.00126827f
cc_24 N_A2_4 N_A3_4 0.00473219f
cc_25 N_MM4_g N_MM5_g 0.00712461f
x_PM_AO33x2_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_AO33x2_ASAP7_75t_R%noxref_16
cc_26 N_noxref_16_1 N_MM24_g 0.00150323f
cc_27 N_noxref_16_1 N_Y_7 0.00074055f
x_PM_AO33x2_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_AO33x2_ASAP7_75t_R%noxref_19
cc_28 N_noxref_19_1 N_NET020_5 0.000502942f
cc_29 N_noxref_19_1 N_NET020_16 0.0345914f
cc_30 N_noxref_19_1 N_MM6_g 0.00233642f
cc_31 N_noxref_19_1 N_noxref_18_1 0.00180995f
x_PM_AO33x2_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_AO33x2_ASAP7_75t_R%noxref_18
cc_32 N_noxref_18_1 N_NET020_16 0.00117077f
cc_33 N_noxref_18_1 N_MM6_g 0.00150044f
x_PM_AO33x2_ASAP7_75t_R%A3 VSS A3 N_MM5_g N_A3_4 N_A3_1 PM_AO33x2_ASAP7_75t_R%A3
cc_34 N_A3_4 N_NET020_1 0.000965285f
cc_35 N_A3_4 N_NET020_19 0.00104114f
cc_36 N_A3_4 N_NET020_18 0.00241054f
cc_37 N_MM5_g N_MM24@2_g 0.00343222f
cc_38 N_A3_4 N_NET020_23 0.00727089f
x_PM_AO33x2_ASAP7_75t_R%Y VSS Y N_MM24_d N_MM24@2_d N_MM25_d N_MM25@2_d N_Y_7
+ N_Y_8 N_Y_9 N_Y_2 N_Y_1 N_Y_14 PM_AO33x2_ASAP7_75t_R%Y
cc_39 N_Y_7 N_NET020_23 0.000209556f
cc_40 N_Y_7 N_NET020_18 0.000339629f
cc_41 N_Y_7 N_NET020_17 0.00124064f
cc_42 N_Y_7 N_NET020_22 0.000451146f
cc_43 N_Y_7 N_NET020_1 0.00538877f
cc_44 N_Y_8 N_MM24@2_g 0.0308453f
cc_45 N_Y_9 N_NET020_17 0.00146084f
cc_46 N_Y_2 N_MM24@2_g 0.00210869f
cc_47 N_Y_1 N_MM24@2_g 0.0022857f
cc_48 N_Y_14 N_NET020_17 0.00251626f
cc_49 N_Y_14 N_NET020_18 0.0033219f
cc_50 N_Y_7 N_MM24_g 0.037088f
cc_51 N_Y_7 N_MM24@2_g 0.0683076f
x_PM_AO33x2_ASAP7_75t_R%B1 VSS B1 N_MM2_g N_B1_1 N_B1_4 PM_AO33x2_ASAP7_75t_R%B1
cc_52 N_MM2_g N_NET020_15 0.0149518f
cc_53 N_B1_1 N_NET020_4 0.000515945f
cc_54 N_B1_4 N_NET020_20 0.000634556f
cc_55 N_MM2_g N_NET020_4 0.00092435f
cc_56 N_B1_4 N_NET020_19 0.00134747f
cc_57 N_B1_1 N_NET020_15 0.00152997f
cc_58 N_MM2_g N_NET020_3 0.00153377f
cc_59 N_B1_4 N_NET020_3 0.00270353f
cc_60 N_MM2_g N_NET020_14 0.0529345f
cc_61 N_B1_4 N_A1_4 0.00361099f
cc_62 N_MM2_g N_MM21_g 0.00594629f
x_PM_AO33x2_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_AO33x2_ASAP7_75t_R%noxref_17
cc_63 N_noxref_17_1 N_MM24_g 0.00149604f
cc_64 N_noxref_17_1 N_Y_8 0.000838122f
cc_65 N_noxref_17_1 N_noxref_16_1 0.00177709f
x_PM_AO33x2_ASAP7_75t_R%B3 VSS B3 N_MM6_g N_B3_1 N_B3_4 PM_AO33x2_ASAP7_75t_R%B3
cc_66 N_MM6_g N_NET020_5 0.00162491f
cc_67 N_B3_1 N_NET020_16 0.000962237f
cc_68 N_B3_4 N_NET020_20 0.00112295f
cc_69 N_B3_4 N_NET020_19 0.00126702f
cc_70 N_B3_4 N_NET020_21 0.00642145f
cc_71 N_MM6_g N_NET020_16 0.0326683f
cc_72 N_B3_1 N_B2_1 0.0013299f
cc_73 N_B3_4 N_B2_4 0.00360567f
cc_74 N_MM6_g N_MM3_g 0.00714858f
x_PM_AO33x2_ASAP7_75t_R%B2 VSS B2 N_MM3_g N_B2_1 N_B2_4 PM_AO33x2_ASAP7_75t_R%B2
cc_75 N_MM3_g N_NET020_3 0.000274399f
cc_76 N_B2_1 N_NET020_4 0.000413971f
cc_77 N_B2_1 N_NET020_15 0.000865077f
cc_78 N_MM3_g N_NET020_4 0.000928339f
cc_79 N_B2_4 N_NET020_20 0.00117901f
cc_80 N_B2_4 N_NET020_19 0.00142443f
cc_81 N_B2_4 N_NET020_4 0.00269443f
cc_82 N_MM3_g N_NET020_15 0.0330702f
cc_83 N_B2_1 N_B1_1 0.00130037f
cc_84 N_B2_4 N_B1_4 0.00335702f
cc_85 N_MM3_g N_MM2_g 0.0070155f
x_PM_AO33x2_ASAP7_75t_R%NET15 VSS N_MM5_d N_MM4_d N_MM21_d N_MM2_s N_MM3_s
+ N_MM6_s N_NET15_13 N_NET15_11 N_NET15_3 N_NET15_12 N_NET15_2 N_NET15_1
+ N_NET15_10 PM_AO33x2_ASAP7_75t_R%NET15
cc_86 N_NET15_13 N_NET020_21 7.45033e-20
cc_87 N_NET15_13 N_NET020_5 0.000206683f
cc_88 N_NET15_13 N_NET020_4 0.000962255f
cc_89 N_NET15_13 N_NET020_16 0.000565729f
cc_90 N_NET15_11 N_NET020_15 0.000603447f
cc_91 N_NET15_3 N_NET020_20 0.00071465f
cc_92 N_NET15_12 N_NET020_15 0.0011346f
cc_93 N_NET15_12 N_NET020_16 0.00113795f
cc_94 N_NET15_2 N_NET020_4 0.00137973f
cc_95 N_NET15_3 N_NET020_4 0.00280153f
cc_96 N_NET15_3 N_NET020_5 0.00442322f
cc_97 N_NET15_13 N_NET020_20 0.0100642f
cc_98 N_NET15_1 N_A3_4 0.00117163f
cc_99 N_NET15_1 N_MM5_g 0.00119674f
cc_100 N_NET15_10 N_MM5_g 0.0329506f
cc_101 N_NET15_10 N_A2_1 0.000661409f
cc_102 N_NET15_13 N_A2_4 0.00115253f
cc_103 N_NET15_1 N_MM4_g 0.00118666f
cc_104 N_NET15_1 N_A2_4 0.00156231f
cc_105 N_NET15_10 N_MM4_g 0.0317493f
cc_106 N_NET15_2 N_MM21_g 0.00118865f
cc_107 N_NET15_13 N_A1_4 0.00123854f
cc_108 N_NET15_2 N_A1_4 0.00176201f
cc_109 N_NET15_11 N_MM21_g 0.0324132f
cc_110 N_NET15_11 N_B1_1 0.000702647f
cc_111 N_NET15_2 N_MM2_g 0.000942193f
cc_112 N_NET15_11 N_MM2_g 0.0321643f
cc_113 N_NET15_12 N_B2_1 0.000696801f
cc_114 N_NET15_3 N_MM3_g 0.000927786f
cc_115 N_NET15_12 N_MM3_g 0.0319744f
cc_116 N_NET15_12 N_B3_1 0.000672631f
cc_117 N_NET15_3 N_MM6_g 0.000928863f
cc_118 N_NET15_12 N_MM6_g 0.0318372f
x_PM_AO33x2_ASAP7_75t_R%NET020 VSS N_MM24_g N_MM24@2_g N_MM7_d N_MM10_d N_MM6_d
+ N_MM2_d N_MM3_d N_NET020_1 N_NET020_19 N_NET020_18 N_NET020_23 N_NET020_14
+ N_NET020_3 N_NET020_20 N_NET020_15 N_NET020_4 N_NET020_5 N_NET020_16
+ N_NET020_21 N_NET020_17 N_NET020_22 PM_AO33x2_ASAP7_75t_R%NET020
*END of AO33x2_ASAP7_75t_R.pxi
.ENDS
** Design:	AOI211x1_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AOI211x1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AOI211x1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AOI211x1_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.0416676f
.ends

.subckt PM_AOI211x1_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.00606965f
.ends

.subckt PM_AOI211x1_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.0420582f
.ends

.subckt PM_AOI211x1_ASAP7_75t_R%NET32 VSS 2 3 1
c1 1 VSS 0.000894844f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_AOI211x1_ASAP7_75t_R%NET17 VSS 19 22 32 35 42 45 10 1 11 2 13 3 12 15
c1 1 VSS 0.00977834f
c2 2 VSS 0.0094796f
c3 3 VSS 0.00330667f
c4 10 VSS 0.00450837f
c5 11 VSS 0.00465501f
c6 12 VSS 0.00236834f
c7 13 VSS 0.0194446f
c8 14 VSS 0.000883589f
c9 15 VSS 0.00330489f
c10 16 VSS 0.000990425f
c11 17 VSS 0.00293291f
r1 45 44 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r2 3 44 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4340 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r3 41 3 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4220 $Y=0.2025 $X2=0.4340 $Y2=0.2025
r4 12 41 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4220 $Y2=0.2025
r5 42 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r6 3 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.1980
r7 37 38 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4095
+ $Y=0.1980 $X2=0.4320 $Y2=0.1980
r8 36 37 7.22888 $w=1.3e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3785
+ $Y=0.1980 $X2=0.4095 $Y2=0.1980
r9 15 16 6.86231 $w=1.42329e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3335 $Y=0.1980 $X2=0.2970 $Y2=0.1980
r10 15 36 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3335
+ $Y=0.1980 $X2=0.3785 $Y2=0.1980
r11 14 17 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.2160 $X2=0.2970 $Y2=0.2340
r12 14 16 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.2160 $X2=0.2970 $Y2=0.1980
r13 35 34 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r14 33 34 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2260 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r15 2 33 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2140 $Y=0.2025 $X2=0.2260 $Y2=0.2025
r16 11 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2140 $Y2=0.2025
r17 32 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r18 17 30 7.32869 $w=1.41688e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.2340 $X2=0.2585 $Y2=0.2340
r19 2 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2150 $Y2=0.2340
r20 29 30 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2270
+ $Y=0.2340 $X2=0.2585 $Y2=0.2340
r21 28 29 0.699569 $w=1.3e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.2240
+ $Y=0.2340 $X2=0.2270 $Y2=0.2340
r22 27 28 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2150
+ $Y=0.2340 $X2=0.2240 $Y2=0.2340
r23 26 27 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1935
+ $Y=0.2340 $X2=0.2150 $Y2=0.2340
r24 25 26 9.79397 $w=1.3e-08 $l=4.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1515
+ $Y=0.2340 $X2=0.1935 $Y2=0.2340
r25 24 25 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1200
+ $Y=0.2340 $X2=0.1515 $Y2=0.2340
r26 23 24 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.1200 $Y2=0.2340
r27 13 23 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.0950
+ $Y=0.2340 $X2=0.1080 $Y2=0.2340
r28 1 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.2340
r29 22 21 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r30 1 21 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1100 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r31 18 1 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0980 $Y=0.2025 $X2=0.1100 $Y2=0.2025
r32 10 18 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.0980 $Y2=0.2025
r33 19 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
.ends

.subckt PM_AOI211x1_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.00537414f
.ends

.subckt PM_AOI211x1_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.0051812f
.ends

.subckt PM_AOI211x1_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.0050782f
.ends

.subckt PM_AOI211x1_ASAP7_75t_R%A1 VSS 23 3 4 8 1 6 9 7
c1 1 VSS 0.0122598f
c2 3 VSS 0.0832698f
c3 4 VSS 0.0844043f
c4 5 VSS 0.00263774f
c5 6 VSS 0.00257868f
c6 7 VSS 0.00332759f
c7 8 VSS 0.0025673f
c8 9 VSS 0.00283879f
r1 9 26 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1980 $X2=0.1890 $Y2=0.1800
r2 25 26 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1620 $X2=0.1890 $Y2=0.1800
r3 6 19 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1485 $X2=0.1890 $Y2=0.1350
r4 6 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1485 $X2=0.1890 $Y2=0.1620
r5 23 24 0.874462 $w=1.3e-08 $l=3.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1190 $X2=0.1890 $Y2=0.1227
r6 23 5 4.4889 $w=1.3e-08 $l=1.93e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1190 $X2=0.1890 $Y2=0.0997
r7 5 7 5.29071 $w=1.46216e-08 $l=2.77e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0997 $X2=0.1890 $Y2=0.0720
r8 4 16 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r9 19 24 1.67627 $w=1.66735e-08 $l=1.23e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1890 $Y2=0.1227
r10 8 18 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2020
+ $Y=0.1350 $X2=0.2130 $Y2=0.1350
r11 8 19 1.85116 $w=1.64615e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2020 $Y=0.1350 $X2=0.1890 $Y2=0.1350
r12 14 16 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2305 $Y=0.1350 $X2=0.2430 $Y2=0.1350
r13 13 14 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2160 $Y=0.1350 $X2=0.2305 $Y2=0.1350
r14 13 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2160 $Y=0.1350
+ $X2=0.2130 $Y2=0.1350
r15 12 13 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2015 $Y=0.1350 $X2=0.2160 $Y2=0.1350
r16 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r17 1 11 3.20232 $w=2.13909e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1780 $Y2=0.1350
r18 1 12 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1890 $Y=0.1350 $X2=0.2015 $Y2=0.1350
r19 3 11 0.905388 $w=2.07755e-07 $l=1.1e-08 $layer=LIG $thickness=5.52727e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1780 $Y2=0.1350
r20 3 12 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1890 $Y=0.1350 $X2=0.2015 $Y2=0.1350
.ends

.subckt PM_AOI211x1_ASAP7_75t_R%B VSS 19 3 4 1 7 6
c1 1 VSS 0.0127578f
c2 3 VSS 0.0478435f
c3 4 VSS 0.045846f
c4 5 VSS 0.00516088f
c5 6 VSS 0.00551806f
c6 7 VSS 0.00416696f
r1 7 21 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.1620 $X2=0.4050 $Y2=0.1485
r2 6 18 4.59114 $w=1.48182e-08 $l=2.47e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.0720 $X2=0.4050 $Y2=0.0967
r3 19 20 1.57403 $w=1.3e-08 $l=6.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1130 $X2=0.4050 $Y2=0.1197
r4 19 18 3.78933 $w=1.3e-08 $l=1.63e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1130 $X2=0.4050 $Y2=0.0967
r5 5 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
r6 5 20 3.55614 $w=1.3e-08 $l=1.53e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1197
r7 5 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1485
r8 3 14 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r9 14 15 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4145 $Y2=0.1350
r10 11 15 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.4175 $Y=0.1350 $X2=0.4145 $Y2=0.1350
r11 10 11 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4320 $Y=0.1350 $X2=0.4175 $Y2=0.1350
r12 9 10 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4465 $Y=0.1350 $X2=0.4320 $Y2=0.1350
r13 4 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r14 1 9 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4465 $Y2=0.1350
r15 1 17 2.90696 $w=2.1681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4695 $Y2=0.1350
r16 4 9 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4465 $Y2=0.1350
r17 4 17 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.4590 $Y=0.1350 $X2=0.4695 $Y2=0.1350
.ends

.subckt PM_AOI211x1_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00552773f
.ends

.subckt PM_AOI211x1_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.00558646f
.ends

.subckt PM_AOI211x1_ASAP7_75t_R%C VSS 25 3 4 1 7 8 6
c1 1 VSS 0.0113544f
c2 3 VSS 0.0451586f
c3 4 VSS 0.0467721f
c4 5 VSS 0.00376507f
c5 6 VSS 0.00465894f
c6 7 VSS 0.0035039f
c7 8 VSS 0.00334132f
r1 25 26 0.524677 $w=1.3e-08 $l=2.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1220 $X2=0.5130 $Y2=0.1242
r2 25 5 4.83869 $w=1.3e-08 $l=2.08e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1220 $X2=0.5130 $Y2=0.1012
r3 5 6 5.64049 $w=1.45385e-08 $l=2.92e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1012 $X2=0.5130 $Y2=0.0720
r4 7 8 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5265 $Y2=0.1350
r5 7 26 1.32648 $w=1.7186e-08 $l=1.08e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5130 $Y2=0.1242
r6 4 17 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1350
r7 8 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5265
+ $Y=0.1350 $X2=0.5400 $Y2=0.1350
r8 15 17 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5545 $Y=0.1350 $X2=0.5670 $Y2=0.1350
r9 14 15 2.36289 $w=1.53e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08 $X=0.5505
+ $Y=0.1350 $X2=0.5545 $Y2=0.1350
r10 13 14 6.20259 $w=1.53e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5400 $Y=0.1350 $X2=0.5505 $Y2=0.1350
r11 13 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5400 $Y=0.1350
+ $X2=0.5400 $Y2=0.1350
r12 12 13 6.20259 $w=1.53e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5295 $Y=0.1350 $X2=0.5400 $Y2=0.1350
r13 11 12 2.36289 $w=1.53e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08 $X=0.5255
+ $Y=0.1350 $X2=0.5295 $Y2=0.1350
r14 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r15 1 10 3.20232 $w=2.13909e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5020 $Y2=0.1350
r16 1 11 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5255 $Y2=0.1350
r17 3 10 0.905388 $w=2.07755e-07 $l=1.1e-08 $layer=LIG $thickness=5.52727e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5020 $Y2=0.1350
r18 3 11 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5255 $Y2=0.1350
.ends

.subckt PM_AOI211x1_ASAP7_75t_R%A2 VSS 25 3 4 1
c1 1 VSS 0.00427525f
c2 3 VSS 0.0436741f
c3 4 VSS 0.0435021f
c4 5 VSS 0.014206f
c5 6 VSS 0.0154835f
c6 7 VSS 0.00514998f
c7 8 VSS 0.00277323f
r1 25 6 1.10765 $w=1.3e-08 $l=4.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1530 $X2=0.0270 $Y2=0.1482
r2 6 8 1.90946 $w=1.63962e-08 $l=1.32e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1482 $X2=0.0270 $Y2=0.1350
r3 5 8 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1035 $X2=0.0270 $Y2=0.1350
r4 8 21 7.33112 $w=1.42329e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1350 $X2=0.0635 $Y2=0.1350
r5 3 16 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r6 7 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0955
+ $Y=0.1350 $X2=0.1090 $Y2=0.1350
r7 7 21 7.46207 $w=1.3e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0955
+ $Y=0.1350 $X2=0.0635 $Y2=0.1350
r8 14 16 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1350 $X2=0.0810 $Y2=0.1350
r9 12 13 5.90723 $w=1.53e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.1090
+ $Y=0.1350 $X2=0.1190 $Y2=0.1350
r10 12 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1090 $Y=0.1350
+ $X2=0.1090 $Y2=0.1350
r11 11 12 6.49795 $w=1.53e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0980 $Y=0.1350 $X2=0.1090 $Y2=0.1350
r12 11 14 2.65825 $w=1.53e-08 $l=4.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0980 $Y=0.1350 $X2=0.0935 $Y2=0.1350
r13 10 13 2.06753 $w=1.53e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1350 $X2=0.1190 $Y2=0.1350
r14 4 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r15 1 10 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1225 $Y2=0.1350
r16 1 18 2.90696 $w=2.1681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1455 $Y2=0.1350
r17 4 10 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1225 $Y2=0.1350
r18 4 18 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.1350 $Y=0.1350 $X2=0.1455 $Y2=0.1350
.ends

.subckt PM_AOI211x1_ASAP7_75t_R%NET34 VSS 16 17 28 30 13 2 1 10 11 3 12
c1 1 VSS 0.00535114f
c2 2 VSS 0.00445185f
c3 3 VSS 0.00541748f
c4 10 VSS 0.00257887f
c5 11 VSS 0.00213184f
c6 12 VSS 0.00233815f
c7 13 VSS 0.0221918f
r1 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2025 $X2=0.5920 $Y2=0.2025
r2 30 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.2025 $X2=0.5795 $Y2=0.2025
r3 28 27 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r4 10 27 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3800 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r5 3 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2025
+ $X2=0.5940 $Y2=0.2340
r6 1 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.2340
r7 24 25 9.79397 $w=1.3e-08 $l=4.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.5520
+ $Y=0.2340 $X2=0.5940 $Y2=0.2340
r8 23 24 9.44418 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.5115
+ $Y=0.2340 $X2=0.5520 $Y2=0.2340
r9 21 22 9.32759 $w=1.3e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.4180 $Y2=0.2340
r10 19 23 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4995
+ $Y=0.2340 $X2=0.5115 $Y2=0.2340
r11 18 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.2340 $X2=0.4995 $Y2=0.2340
r12 13 18 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.4630
+ $Y=0.2340 $X2=0.4860 $Y2=0.2340
r13 13 22 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4630
+ $Y=0.2340 $X2=0.4180 $Y2=0.2340
r14 2 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2025
+ $X2=0.4860 $Y2=0.2340
r15 16 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r16 2 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r17 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4860 $Y2=0.2025
r18 17 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r19 1 10 1e-05
.ends

.subckt PM_AOI211x1_ASAP7_75t_R%Y VSS 40 19 37 38 53 56 1 13 10 11 2 3 12 14 15
+ 17
c1 1 VSS 0.00625134f
c2 2 VSS 0.00996208f
c3 3 VSS 0.00287595f
c4 10 VSS 0.00276238f
c5 11 VSS 0.00452883f
c6 12 VSS 0.00214385f
c7 13 VSS 0.0513508f
c8 14 VSS 0.00118353f
c9 15 VSS 0.00287199f
c10 16 VSS 0.00308827f
c11 17 VSS 0.000773908f
r1 56 55 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r2 54 55 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5500 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r3 3 54 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5380 $Y=0.2025 $X2=0.5500 $Y2=0.2025
r4 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.2025 $X2=0.5380 $Y2=0.2025
r5 53 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.2025 $X2=0.5255 $Y2=0.2025
r6 3 49 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.2025
+ $X2=0.5400 $Y2=0.1980
r7 49 50 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1980 $X2=0.5515 $Y2=0.1980
r8 47 50 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.5810
+ $Y=0.1980 $X2=0.5515 $Y2=0.1980
r9 14 17 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6100 $Y=0.1980 $X2=0.6210 $Y2=0.1980
r10 14 47 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6100
+ $Y=0.1980 $X2=0.5810 $Y2=0.1980
r11 17 46 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1980 $X2=0.6210 $Y2=0.1800
r12 45 46 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1675 $X2=0.6210 $Y2=0.1800
r13 44 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1540 $X2=0.6210 $Y2=0.1675
r14 43 44 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1540
r15 42 43 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1035 $X2=0.6210 $Y2=0.1350
r16 41 42 6.70421 $w=1.3e-08 $l=2.88e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0747 $X2=0.6210 $Y2=0.1035
r17 40 41 1.57403 $w=1.3e-08 $l=6.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0680 $X2=0.6210 $Y2=0.0747
r18 40 39 0.641272 $w=1.3e-08 $l=2.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0680 $X2=0.6210 $Y2=0.0652
r19 15 16 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0540 $X2=0.6210 $Y2=0.0360
r20 15 39 2.62338 $w=1.3e-08 $l=1.12e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0540 $X2=0.6210 $Y2=0.0652
r21 38 36 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0675 $X2=0.5005 $Y2=0.0675
r22 2 36 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.0675 $X2=0.5005 $Y2=0.0675
r23 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0675 $X2=0.4860 $Y2=0.0675
r24 37 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4715 $Y2=0.0675
r25 16 34 7.2121 $w=1.41842e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.0360 $X2=0.5830 $Y2=0.0360
r26 2 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0675
+ $X2=0.4860 $Y2=0.0360
r27 33 34 7.22888 $w=1.3e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5520
+ $Y=0.0360 $X2=0.5830 $Y2=0.0360
r28 32 33 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.5270
+ $Y=0.0360 $X2=0.5520 $Y2=0.0360
r29 31 32 6.41272 $w=1.3e-08 $l=2.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.4995
+ $Y=0.0360 $X2=0.5270 $Y2=0.0360
r30 30 31 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.0360 $X2=0.4995 $Y2=0.0360
r31 29 30 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.4630
+ $Y=0.0360 $X2=0.4860 $Y2=0.0360
r32 28 29 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.4455
+ $Y=0.0360 $X2=0.4630 $Y2=0.0360
r33 27 28 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.4190
+ $Y=0.0360 $X2=0.4455 $Y2=0.0360
r34 26 27 17.9556 $w=1.3e-08 $l=7.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3420
+ $Y=0.0360 $X2=0.4190 $Y2=0.0360
r35 25 26 19.4713 $w=1.3e-08 $l=8.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2585
+ $Y=0.0360 $X2=0.3420 $Y2=0.0360
r36 24 25 7.92845 $w=1.3e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2245
+ $Y=0.0360 $X2=0.2585 $Y2=0.0360
r37 23 24 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.2000
+ $Y=0.0360 $X2=0.2245 $Y2=0.0360
r38 22 23 11.3097 $w=1.3e-08 $l=4.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1515
+ $Y=0.0360 $X2=0.2000 $Y2=0.0360
r39 21 22 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1200
+ $Y=0.0360 $X2=0.1515 $Y2=0.0360
r40 20 21 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.1200 $Y2=0.0360
r41 13 20 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.0950
+ $Y=0.0360 $X2=0.1080 $Y2=0.0360
r42 1 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1080 $Y2=0.0360
r43 19 18 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r44 10 18 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1100 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r45 1 10 1e-05
.ends


*
.SUBCKT AOI211x1_ASAP7_75t_R VSS VDD A2 A1 B C Y
*
* VSS VSS
* VDD VDD
* A2 A2
* A1 A1
* B B
* C C
* Y Y
*
*

MM4 N_MM4_d N_MM4_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM20 N_MM20_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM21 N_MM21_d N_MM21_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM21@2 N_MM21@2_d N_MM4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM5_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@2 N_MM0@2_d N_MM0@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM6_g N_MM6_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6@2 N_MM6@2_d N_MM3_g N_MM6@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM7_g N_MM7_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7@2 N_MM7@2_d N_MM7@2_g N_MM7@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AOI211x1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AOI211x1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AOI211x1_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_AOI211x1_ASAP7_75t_R%noxref_14
cc_1 N_noxref_14_1 N_MM0@2_g 0.00155831f
cc_2 N_noxref_14_1 N_NET34_10 0.000538311f
cc_3 N_noxref_14_1 N_noxref_13_1 0.00138734f
x_PM_AOI211x1_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_AOI211x1_ASAP7_75t_R%noxref_16
cc_4 N_noxref_16_1 N_MM6_g 0.00160108f
cc_5 N_noxref_16_1 N_NET34_10 0.0361613f
cc_6 N_noxref_16_1 N_noxref_13_1 0.000486437f
cc_7 N_noxref_16_1 N_noxref_14_1 0.00766557f
cc_8 N_noxref_16_1 N_noxref_15_1 0.00138037f
x_PM_AOI211x1_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_AOI211x1_ASAP7_75t_R%noxref_12
cc_9 N_noxref_12_1 N_MM21_g 0.00247486f
cc_10 N_noxref_12_1 N_noxref_11_1 0.00194752f
x_PM_AOI211x1_ASAP7_75t_R%NET32 VSS N_MM4_s N_MM5_d N_NET32_1
+ PM_AOI211x1_ASAP7_75t_R%NET32
cc_11 N_NET32_1 N_MM4_g 0.0172615f
cc_12 N_NET32_1 N_MM5_g 0.0172889f
x_PM_AOI211x1_ASAP7_75t_R%NET17 VSS N_MM21_d N_MM21@2_d N_MM0_d N_MM0@2_d
+ N_MM6_s N_MM6@2_s N_NET17_10 N_NET17_1 N_NET17_11 N_NET17_2 N_NET17_13
+ N_NET17_3 N_NET17_12 N_NET17_15 PM_AOI211x1_ASAP7_75t_R%NET17
cc_13 N_NET17_10 N_A2_1 0.0020571f
cc_14 N_NET17_1 N_MM4_g 0.0021645f
cc_15 N_NET17_10 N_MM21_g 0.0181454f
cc_16 N_NET17_10 N_MM4_g 0.050788f
cc_17 N_NET17_11 N_A1_6 0.000641718f
cc_18 N_NET17_11 N_A1_1 0.0020348f
cc_19 N_NET17_2 N_MM0@2_g 0.00249834f
cc_20 N_NET17_13 N_A1_9 0.00571284f
cc_21 N_NET17_11 N_MM5_g 0.0181691f
cc_22 N_NET17_11 N_MM0@2_g 0.050294f
cc_23 N_NET17_3 N_MM3_g 0.00198924f
cc_24 N_NET17_12 N_B_1 0.00210713f
cc_25 N_NET17_15 N_B_7 0.00527633f
cc_26 N_NET17_12 N_MM6_g 0.0181888f
cc_27 N_NET17_12 N_MM3_g 0.0495243f
x_PM_AOI211x1_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_AOI211x1_ASAP7_75t_R%noxref_11
cc_28 N_noxref_11_1 N_MM21_g 0.010424f
cc_29 N_noxref_11_1 N_Y_10 0.000632695f
x_PM_AOI211x1_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_AOI211x1_ASAP7_75t_R%noxref_17
cc_30 N_noxref_17_1 N_MM7@2_g 0.00916427f
cc_31 N_noxref_17_1 N_NET34_12 0.000631095f
cc_32 N_noxref_17_1 N_Y_15 0.00136337f
x_PM_AOI211x1_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_AOI211x1_ASAP7_75t_R%noxref_15
cc_33 N_noxref_15_1 N_MM0@2_g 0.000288518f
cc_34 N_noxref_15_1 N_MM6_g 0.00924482f
cc_35 N_noxref_15_1 N_NET34_10 0.000527504f
cc_36 N_noxref_15_1 N_Y_13 0.000519828f
cc_37 N_noxref_15_1 N_noxref_13_1 0.00804513f
cc_38 N_noxref_15_1 N_noxref_14_1 0.00048362f
x_PM_AOI211x1_ASAP7_75t_R%A1 VSS A1 N_MM5_g N_MM0@2_g N_A1_8 N_A1_1 N_A1_6
+ N_A1_9 N_A1_7 PM_AOI211x1_ASAP7_75t_R%A1
cc_39 N_A1_8 N_MM4_g 0.000902931f
cc_40 N_A1_1 N_A2_1 0.00150127f
cc_41 N_MM5_g N_MM4_g 0.00664578f
x_PM_AOI211x1_ASAP7_75t_R%B VSS B N_MM6_g N_MM3_g N_B_1 N_B_7 N_B_6
+ PM_AOI211x1_ASAP7_75t_R%B
x_PM_AOI211x1_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_AOI211x1_ASAP7_75t_R%noxref_13
cc_42 N_noxref_13_1 N_MM0@2_g 0.00909182f
cc_43 N_noxref_13_1 N_MM6_g 0.000490404f
cc_44 N_noxref_13_1 N_Y_13 0.000540237f
x_PM_AOI211x1_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_AOI211x1_ASAP7_75t_R%noxref_18
cc_45 N_noxref_18_1 N_MM7@2_g 0.00164206f
cc_46 N_noxref_18_1 N_NET34_12 0.036501f
cc_47 N_noxref_18_1 N_Y_12 0.000778436f
cc_48 N_noxref_18_1 N_noxref_17_1 0.00193956f
x_PM_AOI211x1_ASAP7_75t_R%C VSS C N_MM7_g N_MM7@2_g N_C_1 N_C_7 N_C_8 N_C_6
+ PM_AOI211x1_ASAP7_75t_R%C
cc_49 N_MM7_g N_B_1 0.0012399f
cc_50 N_MM7_g N_MM3_g 0.00534403f
x_PM_AOI211x1_ASAP7_75t_R%A2 VSS A2 N_MM21_g N_MM4_g N_A2_1
+ PM_AOI211x1_ASAP7_75t_R%A2
x_PM_AOI211x1_ASAP7_75t_R%NET34 VSS N_MM7_s N_MM6@2_d N_MM6_d N_MM7@2_s
+ N_NET34_13 N_NET34_2 N_NET34_1 N_NET34_10 N_NET34_11 N_NET34_3 N_NET34_12
+ PM_AOI211x1_ASAP7_75t_R%NET34
cc_51 N_NET34_13 N_MM6_g 0.000503856f
cc_52 N_NET34_2 N_MM3_g 0.000833011f
cc_53 N_NET34_1 N_MM6_g 0.00121988f
cc_54 N_NET34_10 N_B_1 0.00160407f
cc_55 N_NET34_11 N_MM3_g 0.0333385f
cc_56 N_NET34_10 N_MM6_g 0.0354209f
cc_57 N_NET34_11 N_MM7@2_g 0.000469927f
cc_58 N_NET34_2 N_MM7@2_g 0.000980529f
cc_59 N_NET34_3 N_MM7@2_g 0.00103315f
cc_60 N_NET34_12 N_C_1 0.0017687f
cc_61 N_NET34_11 N_MM7_g 0.0334427f
cc_62 N_NET34_12 N_MM7@2_g 0.0353902f
cc_63 N_NET34_10 N_NET17_15 0.000625509f
cc_64 N_NET34_1 N_NET17_15 0.000627185f
cc_65 N_NET34_11 N_NET17_12 0.00110753f
cc_66 N_NET34_1 N_NET17_3 0.00211201f
cc_67 N_NET34_2 N_NET17_3 0.00415011f
cc_68 N_NET34_13 N_NET17_15 0.0111967f
x_PM_AOI211x1_ASAP7_75t_R%Y VSS Y N_MM4_d N_MM3_d N_MM20_d N_MM7_d N_MM7@2_d
+ N_Y_1 N_Y_13 N_Y_10 N_Y_11 N_Y_2 N_Y_3 N_Y_12 N_Y_14 N_Y_15 N_Y_17
+ PM_AOI211x1_ASAP7_75t_R%Y
cc_69 N_Y_1 N_MM4_g 0.00368297f
cc_70 N_Y_13 N_MM4_g 0.00158248f
cc_71 N_Y_10 N_A2_1 0.00235146f
cc_72 N_Y_10 N_MM21_g 0.019056f
cc_73 N_Y_10 N_MM4_g 0.0531829f
cc_74 N_Y_10 N_A1_7 0.000261553f
cc_75 N_Y_1 N_A1_7 0.00035354f
cc_76 N_Y_13 N_A1_7 0.007233f
cc_77 N_Y_13 N_MM3_g 0.000597126f
cc_78 N_Y_11 N_B_1 0.000930474f
cc_79 N_Y_2 N_MM3_g 0.000968315f
cc_80 N_Y_13 N_B_6 0.00576426f
cc_81 N_Y_11 N_MM3_g 0.0347065f
cc_82 N_Y_3 N_MM7_g 0.000633685f
cc_83 N_Y_2 N_MM7_g 0.0020641f
cc_84 N_Y_12 N_MM7_g 0.000808373f
cc_85 N_Y_14 N_C_7 0.00104133f
cc_86 N_Y_15 N_C_1 0.00137336f
cc_87 N_Y_3 N_MM7@2_g 0.00196228f
cc_88 N_Y_14 N_C_8 0.00215244f
cc_89 N_Y_12 N_C_1 0.00347689f
cc_90 N_Y_13 N_C_6 0.00596705f
cc_91 N_Y_12 N_MM7@2_g 0.0488484f
cc_92 N_Y_11 N_MM7_g 0.0533224f
cc_93 N_Y_12 N_NET34_13 0.000599342f
cc_94 N_Y_17 N_NET34_13 0.000625995f
cc_95 N_Y_3 N_NET34_13 0.000651013f
cc_96 N_Y_14 N_NET34_3 0.000682429f
cc_97 N_Y_12 N_NET34_12 0.00182069f
cc_98 N_Y_15 N_NET34_3 0.000798809f
cc_99 N_Y_3 N_NET34_2 0.00145569f
cc_100 N_Y_3 N_NET34_3 0.00527351f
cc_101 N_Y_14 N_NET34_13 0.00948633f
*END of AOI211x1_ASAP7_75t_R.pxi
.ENDS
** Design:	AOI211xp5_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AOI211xp5_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AOI211xp5_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AOI211xp5_ASAP7_75t_R%NET34 VSS 2 3 1
c1 1 VSS 0.000978869f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2160 $Y2=0.2025
.ends

.subckt PM_AOI211xp5_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.042167f
.ends

.subckt PM_AOI211xp5_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.0322608f
.ends

.subckt PM_AOI211xp5_ASAP7_75t_R%C VSS 6 3 1 4
c1 1 VSS 0.00495803f
c2 3 VSS 0.0728053f
c3 4 VSS 0.00293218f
r1 7 8 2.39019 $w=1.3e-08 $l=1.03e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1247 $X2=0.2430 $Y2=0.1350
r2 6 7 0.408082 $w=1.3e-08 $l=1.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1230 $X2=0.2430 $Y2=0.1247
r3 6 4 6.23783 $w=1.3e-08 $l=2.68e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1230 $X2=0.2430 $Y2=0.0962
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AOI211xp5_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.00574318f
.ends

.subckt PM_AOI211xp5_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.00459195f
.ends

.subckt PM_AOI211xp5_ASAP7_75t_R%NET32 VSS 2 3 1
c1 1 VSS 0.000861305f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0540 $X2=0.1080 $Y2=0.0540
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0540 $X2=0.1080 $Y2=0.0540
.ends

.subckt PM_AOI211xp5_ASAP7_75t_R%NET17 VSS 11 20 21 7 9 1 8 2
c1 1 VSS 0.00538617f
c2 2 VSS 0.00576291f
c3 7 VSS 0.00221593f
c4 8 VSS 0.0028282f
c5 9 VSS 0.0124807f
r1 21 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r2 2 19 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r4 20 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r5 2 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r6 15 16 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.1260
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r7 14 15 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.2340 $X2=0.1260 $Y2=0.2340
r8 13 14 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0765
+ $Y=0.2340 $X2=0.0945 $Y2=0.2340
r9 12 13 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2340 $X2=0.0765 $Y2=0.2340
r10 9 12 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r11 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r12 11 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r13 7 10 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r14 1 7 1e-05
.ends

.subckt PM_AOI211xp5_ASAP7_75t_R%Y VSS 38 19 34 35 50 51 10 2 12 13 1 14 3 11
+ 15 17
c1 1 VSS 0.00615606f
c2 2 VSS 0.00290305f
c3 3 VSS 0.00841861f
c4 10 VSS 0.00262131f
c5 11 VSS 0.00394309f
c6 12 VSS 0.0022924f
c7 13 VSS 0.0235256f
c8 14 VSS 0.00584847f
c9 15 VSS 0.00480811f
c10 16 VSS 0.00343216f
c11 17 VSS 0.00164634f
r1 51 49 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r2 2 49 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r3 12 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r4 50 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
r5 2 46 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.1980
r6 46 47 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.1980 $X2=0.1215 $Y2=0.1980
r7 45 47 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1980 $X2=0.1215 $Y2=0.1980
r8 44 45 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1600
+ $Y=0.1980 $X2=0.1350 $Y2=0.1980
r9 43 44 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1780
+ $Y=0.1980 $X2=0.1600 $Y2=0.1980
r10 42 43 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1980 $X2=0.1780 $Y2=0.1980
r11 41 42 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1980 $X2=0.1890 $Y2=0.1980
r12 40 41 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1980 $X2=0.2160 $Y2=0.1980
r13 14 17 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2700 $Y=0.1980 $X2=0.2970 $Y2=0.1980
r14 14 40 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1980 $X2=0.2430 $Y2=0.1980
r15 17 39 2.37341 $w=1.8113e-08 $l=1.73e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1980 $X2=0.2970 $Y2=0.1807
r16 38 39 2.04041 $w=1.3e-08 $l=8.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1720 $X2=0.2970 $Y2=0.1807
r17 38 37 0.991056 $w=1.3e-08 $l=4.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1720 $X2=0.2970 $Y2=0.1677
r18 36 37 11.8344 $w=1.3e-08 $l=5.07e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1170 $X2=0.2970 $Y2=0.1677
r19 15 16 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0575 $X2=0.2970 $Y2=0.0360
r20 15 36 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0575 $X2=0.2970 $Y2=0.1170
r21 35 33 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0540 $X2=0.2305 $Y2=0.0540
r22 3 33 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.0540 $X2=0.2305 $Y2=0.0540
r23 11 3 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0540 $X2=0.2160 $Y2=0.0540
r24 34 11 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0540 $X2=0.2015 $Y2=0.0540
r25 16 31 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0360 $X2=0.2700 $Y2=0.0360
r26 3 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0540
+ $X2=0.2160 $Y2=0.0360
r27 30 31 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r28 29 30 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r29 28 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.2295 $Y2=0.0360
r30 27 28 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2025
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r31 26 27 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.2025 $Y2=0.0360
r32 25 26 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r33 24 25 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r34 23 24 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1125
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r35 22 23 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.0360 $X2=0.1125 $Y2=0.0360
r36 21 22 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0765
+ $Y=0.0360 $X2=0.0945 $Y2=0.0360
r37 20 21 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.0360 $X2=0.0765 $Y2=0.0360
r38 13 20 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r39 1 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0540 $Y2=0.0360
r40 19 18 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r41 10 18 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r42 1 10 1e-05
.ends

.subckt PM_AOI211xp5_ASAP7_75t_R%B VSS 8 3 1 4
c1 1 VSS 0.00561151f
c2 3 VSS 0.035214f
c3 4 VSS 0.00377372f
r1 8 7 0.524677 $w=1.3e-08 $l=2.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1480 $X2=0.1890 $Y2=0.1457
r2 6 7 2.50679 $w=1.3e-08 $l=1.07e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1457
r3 4 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0980 $X2=0.1890 $Y2=0.1350
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r5 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AOI211xp5_ASAP7_75t_R%A1 VSS 7 3 1 4
c1 1 VSS 0.00544275f
c2 3 VSS 0.0352809f
c3 4 VSS 0.00393737f
r1 7 8 2.04041 $w=1.3e-08 $l=8.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1090 $X2=0.1350 $Y2=0.1177
r2 4 8 4.02252 $w=1.3e-08 $l=1.73e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1177
r3 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r4 1 4 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AOI211xp5_ASAP7_75t_R%A2 VSS 12 3 1 6 5 4
c1 1 VSS 0.00041191f
c2 3 VSS 0.00533579f
c3 4 VSS 0.00717212f
c4 5 VSS 0.00698407f
c5 6 VSS 0.00251479f
c6 7 VSS 0.00223738f
r1 12 11 2.73998 $w=1.3e-08 $l=1.18e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1870 $X2=0.0270 $Y2=0.1752
r2 5 7 3.2503 $w=1.53684e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1540 $X2=0.0270 $Y2=0.1350
r3 5 11 4.95528 $w=1.3e-08 $l=2.12e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1540 $X2=0.0270 $Y2=0.1752
r4 4 7 7.44771 $w=1.42162e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0980 $X2=0.0270 $Y2=0.1350
r5 7 10 1.38478 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1350 $X2=0.0380 $Y2=0.1350
r6 6 9 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.0560
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r7 6 10 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0560
+ $Y=0.1350 $X2=0.0380 $Y2=0.1350
r8 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r9 1 9 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends


*
.SUBCKT AOI211xp5_ASAP7_75t_R VSS VDD A2 A1 B C Y
*
* VSS VSS
* VDD VDD
* A2 A2
* A1 A1
* B B
* C C
* Y Y
*
*

MM4 N_MM4_d N_MM4_g N_MM4_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM5_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM20 N_MM20_d N_MM20_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM21 N_MM21_d N_MM4_g N_MM21_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM5_g N_MM0_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM3_g N_MM6_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 VDD N_MM20_g N_MM7_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AOI211xp5_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AOI211xp5_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AOI211xp5_ASAP7_75t_R%NET34 VSS N_MM6_d N_MM7_s N_NET34_1
+ PM_AOI211xp5_ASAP7_75t_R%NET34
cc_1 N_NET34_1 N_MM3_g 0.0173175f
cc_2 N_NET34_1 N_MM20_g 0.0174117f
x_PM_AOI211xp5_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_AOI211xp5_ASAP7_75t_R%noxref_14
cc_3 N_noxref_14_1 N_MM20_g 0.00158631f
cc_4 N_noxref_14_1 N_Y_17 0.000736101f
cc_5 N_noxref_14_1 N_noxref_13_1 0.00189611f
x_PM_AOI211xp5_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_AOI211xp5_ASAP7_75t_R%noxref_13
cc_6 N_noxref_13_1 N_MM20_g 0.00348104f
cc_7 N_noxref_13_1 N_Y_11 0.000996657f
x_PM_AOI211xp5_ASAP7_75t_R%C VSS C N_MM20_g N_C_1 N_C_4
+ PM_AOI211xp5_ASAP7_75t_R%C
cc_8 N_C_1 N_B_1 0.00154879f
cc_9 N_C_4 N_B_4 0.00326444f
cc_10 N_MM20_g N_MM3_g 0.00806391f
x_PM_AOI211xp5_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_AOI211xp5_ASAP7_75t_R%noxref_12
cc_11 N_noxref_12_1 N_MM4_g 0.00224272f
cc_12 N_noxref_12_1 N_NET17_7 0.0365376f
cc_13 N_noxref_12_1 N_noxref_11_1 0.00190164f
x_PM_AOI211xp5_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_AOI211xp5_ASAP7_75t_R%noxref_11
cc_14 N_noxref_11_1 N_MM4_g 0.00421035f
cc_15 N_noxref_11_1 N_NET17_7 0.000598308f
cc_16 N_noxref_11_1 N_Y_10 0.0272944f
x_PM_AOI211xp5_ASAP7_75t_R%NET32 VSS N_MM4_s N_MM5_d N_NET32_1
+ PM_AOI211xp5_ASAP7_75t_R%NET32
cc_17 N_NET32_1 N_MM4_g 0.0124889f
cc_18 N_NET32_1 N_MM5_g 0.0125351f
x_PM_AOI211xp5_ASAP7_75t_R%NET17 VSS N_MM21_d N_MM0_d N_MM6_s N_NET17_7
+ N_NET17_9 N_NET17_1 N_NET17_8 N_NET17_2 PM_AOI211xp5_ASAP7_75t_R%NET17
cc_19 N_NET17_7 N_A2_1 0.00066651f
cc_20 N_NET17_9 N_A2_5 0.000901271f
cc_21 N_NET17_1 N_A2_5 0.00147951f
cc_22 N_NET17_1 N_MM4_g 0.00184851f
cc_23 N_NET17_7 N_MM4_g 0.0352739f
cc_24 N_NET17_8 N_A1_1 0.000602315f
cc_25 N_NET17_2 N_MM5_g 0.00092133f
cc_26 N_NET17_8 N_MM5_g 0.0344957f
cc_27 N_NET17_8 N_B_1 0.000857144f
cc_28 N_NET17_2 N_MM3_g 0.00120627f
cc_29 N_NET17_8 N_MM3_g 0.0349358f
x_PM_AOI211xp5_ASAP7_75t_R%Y VSS Y N_MM4_d N_MM3_d N_MM20_d N_MM21_s N_MM0_s
+ N_Y_10 N_Y_2 N_Y_12 N_Y_13 N_Y_1 N_Y_14 N_Y_3 N_Y_11 N_Y_15 N_Y_17
+ PM_AOI211xp5_ASAP7_75t_R%Y
cc_30 N_Y_10 N_MM4_g 0.0112818f
cc_31 N_Y_2 N_A2_1 0.000554763f
cc_32 N_Y_2 N_MM4_g 0.000926509f
cc_33 N_Y_12 N_A2_1 0.0009504f
cc_34 N_Y_13 N_A2_6 0.00113618f
cc_35 N_Y_1 N_MM4_g 0.00123424f
cc_36 N_Y_14 N_A2_6 0.00126063f
cc_37 N_Y_13 N_A2_4 0.00142934f
cc_38 N_Y_12 N_MM4_g 0.0494717f
cc_39 N_Y_12 N_A1_1 0.000751842f
cc_40 N_Y_2 N_MM5_g 0.000921729f
cc_41 N_Y_14 N_A1_4 0.00123992f
cc_42 N_Y_13 N_A1_4 0.00151281f
cc_43 N_Y_2 N_A1_4 0.00287266f
cc_44 N_Y_12 N_MM5_g 0.0358881f
cc_45 N_Y_3 N_MM3_g 0.000665992f
cc_46 N_Y_13 N_B_4 0.00123135f
cc_47 N_Y_14 N_B_4 0.0014464f
cc_48 N_Y_3 N_B_4 0.00283715f
cc_49 N_Y_11 N_MM3_g 0.0258811f
cc_50 N_Y_15 N_C_1 0.000542262f
cc_51 N_Y_3 N_MM20_g 0.000706413f
cc_52 N_Y_13 N_C_4 0.00112349f
cc_53 N_Y_14 N_C_4 0.00138079f
cc_54 N_Y_15 N_C_4 0.00646844f
cc_55 N_Y_11 N_MM20_g 0.0256795f
cc_56 N_Y_12 N_NET17_7 0.000598693f
cc_57 N_Y_12 N_NET17_8 0.00174342f
cc_58 N_Y_2 N_NET17_9 0.000790563f
cc_59 N_Y_2 N_NET17_1 0.00144478f
cc_60 N_Y_2 N_NET17_2 0.00487726f
cc_61 N_Y_14 N_NET17_9 0.0100346f
x_PM_AOI211xp5_ASAP7_75t_R%B VSS B N_MM3_g N_B_1 N_B_4
+ PM_AOI211xp5_ASAP7_75t_R%B
cc_62 N_B_1 N_A1_1 0.00126724f
cc_63 N_B_4 N_A1_4 0.00343016f
cc_64 N_MM3_g N_MM5_g 0.00625103f
x_PM_AOI211xp5_ASAP7_75t_R%A1 VSS A1 N_MM5_g N_A1_1 N_A1_4
+ PM_AOI211xp5_ASAP7_75t_R%A1
cc_65 N_A1_1 N_A2_1 0.00133084f
cc_66 N_A1_4 N_A2_6 0.00201729f
cc_67 N_MM5_g N_MM4_g 0.00789848f
x_PM_AOI211xp5_ASAP7_75t_R%A2 VSS A2 N_MM4_g N_A2_1 N_A2_6 N_A2_5 N_A2_4
+ PM_AOI211xp5_ASAP7_75t_R%A2
*END of AOI211xp5_ASAP7_75t_R.pxi
.ENDS
** Design:	AOI21x1_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AOI21x1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AOI21x1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AOI21x1_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.0315998f
.ends

.subckt PM_AOI21x1_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.0315962f
.ends

.subckt PM_AOI21x1_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.00498956f
.ends

.subckt PM_AOI21x1_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00492295f
.ends

.subckt PM_AOI21x1_ASAP7_75t_R%NET29__2 VSS 2 3 1
c1 1 VSS 0.000962842f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_AOI21x1_ASAP7_75t_R%A2 VSS 5 3 4 1 6
c1 1 VSS 0.0135344f
c2 3 VSS 0.0845297f
c3 4 VSS 0.0846446f
c4 5 VSS 0.00474935f
c5 6 VSS 0.00286763f
r1 5 6 0.763861 $w=3.26364e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2085 $Y=0.1340 $X2=0.2290 $Y2=0.1340
r2 6 18 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2290
+ $Y=0.1340 $X2=0.2400 $Y2=0.1340
r3 4 15 0.314665 $w=2.27e-07 $l=0 $layer=Gate_1 $thickness=5.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r4 13 15 2.08928 $w=2.2e-08 $l=2e-09 $layer=LIG $thickness=4.8e-08 $X=0.2410
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r5 13 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2410 $Y=0.1350
+ $X2=0.2400 $Y2=0.1340
r6 12 13 2.68 $w=2.12556e-08 $l=9e-09 $layer=LIG $thickness=4.8e-08 $X=0.2320
+ $Y=0.1350 $X2=0.2410 $Y2=0.1350
r7 11 12 1.47681 $w=1.53e-08 $l=2.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2295
+ $Y=0.1350 $X2=0.2320 $Y2=0.1350
r8 10 11 7.97476 $w=1.53e-08 $l=1.35e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2160 $Y=0.1350 $X2=0.2295 $Y2=0.1350
r9 9 10 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08 $X=0.2015
+ $Y=0.1350 $X2=0.2160 $Y2=0.1350
r10 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r11 1 8 3.05464 $w=2.15326e-08 $l=1.08e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1782 $Y2=0.1350
r12 1 9 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1890 $Y=0.1350 $X2=0.2015 $Y2=0.1350
r13 3 8 0.757708 $w=2.1223e-07 $l=1.08e-08 $layer=LIG $thickness=5.54419e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1782 $Y2=0.1350
r14 3 9 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1890 $Y=0.1350 $X2=0.2015 $Y2=0.1350
.ends

.subckt PM_AOI21x1_ASAP7_75t_R%NET29 VSS 2 3 1
c1 1 VSS 0.000968907f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2700 $Y2=0.0675
.ends

.subckt PM_AOI21x1_ASAP7_75t_R%NET18 VSS 15 18 24 27 30 31 10 1 2 12 3 13 11
c1 1 VSS 0.00701161f
c2 2 VSS 0.00896286f
c3 3 VSS 0.00685071f
c4 10 VSS 0.00324666f
c5 11 VSS 0.00442764f
c6 12 VSS 0.00324915f
c7 13 VSS 0.0228952f
r1 31 29 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r2 2 29 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r3 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r4 30 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r5 27 26 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r6 1 26 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1100 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r7 23 1 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0980 $Y=0.2025 $X2=0.1100 $Y2=0.2025
r8 10 23 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.0980 $Y2=0.2025
r9 24 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
r10 2 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.2340
r11 1 13 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.2340
r12 21 22 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.3240 $Y2=0.2340
r13 20 21 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r14 19 20 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r15 13 19 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r16 3 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.2340
r17 18 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r18 16 17 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3340 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r19 3 16 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3220 $Y=0.2025 $X2=0.3340 $Y2=0.2025
r20 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3220 $Y2=0.2025
r21 15 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
.ends

.subckt PM_AOI21x1_ASAP7_75t_R%B VSS 15 5 6 2 1 8 9 7 11 10
c1 1 VSS 0.00553844f
c2 2 VSS 0.00547286f
c3 5 VSS 0.0339453f
c4 6 VSS 0.0339583f
c5 7 VSS 0.00364573f
c6 8 VSS 0.00712145f
c7 9 VSS 0.0029738f
c8 10 VSS 0.00262378f
c9 11 VSS 0.00260327f
r1 2 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1340
r2 6 2 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r3 30 31 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1340 $X2=0.3510 $Y2=0.1535
r4 28 31 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1675 $X2=0.3510 $Y2=0.1535
r5 9 11 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1800 $X2=0.3510 $Y2=0.1980
r6 9 28 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1800 $X2=0.3510 $Y2=0.1675
r7 11 27 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.1980 $X2=0.3375 $Y2=0.1980
r8 26 27 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3195
+ $Y=0.1980 $X2=0.3375 $Y2=0.1980
r9 25 26 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1980 $X2=0.3195 $Y2=0.1980
r10 24 25 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2720
+ $Y=0.1980 $X2=0.2970 $Y2=0.1980
r11 23 24 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2415
+ $Y=0.1980 $X2=0.2720 $Y2=0.1980
r12 22 23 7.69526 $w=1.3e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.2085
+ $Y=0.1980 $X2=0.2415 $Y2=0.1980
r13 21 22 9.67737 $w=1.3e-08 $l=4.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1670
+ $Y=0.1980 $X2=0.2085 $Y2=0.1980
r14 20 21 7.46207 $w=1.3e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1980 $X2=0.1670 $Y2=0.1980
r15 19 20 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1125
+ $Y=0.1980 $X2=0.1350 $Y2=0.1980
r16 8 10 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.1980 $X2=0.0810 $Y2=0.1980
r17 8 19 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.1980 $X2=0.1125 $Y2=0.1980
r18 10 18 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1980 $X2=0.0810 $Y2=0.1800
r19 17 18 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1675 $X2=0.0810 $Y2=0.1800
r20 16 17 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1535 $X2=0.0810 $Y2=0.1675
r21 15 16 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1340 $X2=0.0810 $Y2=0.1535
r22 15 7 8.51143 $w=1.3e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1340 $X2=0.0810 $Y2=0.0975
r23 5 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r24 15 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1340
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AOI21x1_ASAP7_75t_R%A1 VSS 24 5 6 7 2 1 9 8 10 11
c1 1 VSS 0.00630455f
c2 2 VSS 0.00633884f
c3 5 VSS 0.0454537f
c4 6 VSS 0.0454686f
c5 7 VSS 0.00310202f
c6 8 VSS 0.00526987f
c7 9 VSS 0.00312113f
c8 10 VSS 0.00241128f
c9 11 VSS 0.00255839f
r1 24 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1340
+ $X2=0.1350 $Y2=0.1350
r2 5 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r3 24 23 5.13017 $w=1.3e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1340 $X2=0.1350 $Y2=0.1120
r4 7 22 2.65995 $w=1.48966e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.0900 $X2=0.1350 $Y2=0.0755
r5 7 23 5.13017 $w=1.3e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0900 $X2=0.1350 $Y2=0.1120
r6 10 21 5.72052 $w=1.36604e-08 $l=3.24692e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.0665 $X2=0.1670 $Y2=0.0720
r7 10 22 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0665 $X2=0.1350 $Y2=0.0755
r8 20 21 9.67737 $w=1.3e-08 $l=4.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2085
+ $Y=0.0720 $X2=0.1670 $Y2=0.0720
r9 19 20 7.69526 $w=1.3e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.2415
+ $Y=0.0720 $X2=0.2085 $Y2=0.0720
r10 8 11 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2720
+ $Y=0.0720 $X2=0.2970 $Y2=0.0720
r11 8 19 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2720
+ $Y=0.0720 $X2=0.2415 $Y2=0.0720
r12 11 17 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0720 $X2=0.2970 $Y2=0.0900
r13 16 17 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1075 $X2=0.2970 $Y2=0.0900
r14 15 16 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1205 $X2=0.2970 $Y2=0.1075
r15 9 15 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1340 $X2=0.2970 $Y2=0.1205
r16 6 2 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r17 2 9 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1340
.ends

.subckt PM_AOI21x1_ASAP7_75t_R%Y VSS 52 30 31 57 58 71 73 1 4 14 16 19 2 3 22
+ 26 25 20 23 21 15 13
c1 1 VSS 0.00531874f
c2 2 VSS 0.00748209f
c3 3 VSS 0.007829f
c4 4 VSS 0.00549886f
c5 13 VSS 0.00335642f
c6 14 VSS 0.000612742f
c7 15 VSS 0.00315267f
c8 16 VSS 0.000613801f
c9 17 VSS 5.68827e-20
c10 18 VSS 5.57833e-20
c11 19 VSS 0.0023724f
c12 20 VSS 0.00237363f
c13 21 VSS 0.00402731f
c14 22 VSS 0.0333711f
c15 23 VSS 0.00433965f
c16 24 VSS 0.0034506f
c17 25 VSS 0.00550292f
c18 26 VSS 0.00461676f
c19 27 VSS 0.0034276f
r1 20 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3760 $Y2=0.2025
r2 73 20 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r3 71 70 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r4 19 70 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r5 4 68 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.2340
r6 1 67 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r7 68 69 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r8 26 65 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.2340 $X2=0.4050 $Y2=0.2160
r9 26 69 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.2340 $X2=0.3915 $Y2=0.2340
r10 66 67 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r11 25 54 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.2340 $X2=0.0270 $Y2=0.2160
r12 25 66 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0405 $Y2=0.2340
r13 64 65 12.7088 $w=1.3e-08 $l=5.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1615 $X2=0.4050 $Y2=0.2160
r14 63 64 16.7897 $w=1.3e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0895 $X2=0.4050 $Y2=0.1615
r15 23 27 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0540 $X2=0.4050 $Y2=0.0360
r16 23 63 8.27824 $w=1.3e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0540 $X2=0.4050 $Y2=0.0895
r17 61 62 0.264706 $w=1.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3340 $Y=0.0725 $X2=0.3385 $Y2=0.0725
r18 3 61 0.705882 $w=1.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3220 $Y=0.0725 $X2=0.3340 $Y2=0.0725
r19 18 3 0.735294 $w=1.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0725 $X2=0.3220 $Y2=0.0725
r20 16 3 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0945 $X2=0.3220 $Y2=0.0945
r21 58 56 0.0675676 $w=3.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0455 $X2=0.3385 $Y2=0.0455
r22 3 56 0.391892 $w=3.7e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.0455 $X2=0.3385 $Y2=0.0455
r23 3 62 0.471383 $w=3.35517e-08 $l=3.06472e-08 $layer=N_src_drn
+ $thickness=1e-09 $X=0.3240 $Y=0.0455 $X2=0.3385 $Y2=0.0725
r24 15 3 0.391892 $w=3.7e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0455 $X2=0.3240 $Y2=0.0455
r25 57 15 0.0675676 $w=3.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0455 $X2=0.3095 $Y2=0.0455
r26 53 54 13.2335 $w=1.3e-08 $l=5.68e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1592 $X2=0.0270 $Y2=0.2160
r27 52 53 11.2514 $w=1.3e-08 $l=4.82e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1110 $X2=0.0270 $Y2=0.1592
r28 52 51 4.83869 $w=1.3e-08 $l=2.08e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1110 $X2=0.0270 $Y2=0.0902
r29 50 51 5.53826 $w=1.3e-08 $l=2.37e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0665 $X2=0.0270 $Y2=0.0902
r30 21 24 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0540 $X2=0.0270 $Y2=0.0360
r31 21 50 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0540 $X2=0.0270 $Y2=0.0665
r32 27 48 3.59766 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0360 $X2=0.3825 $Y2=0.0360
r33 3 44 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0540
+ $X2=0.3240 $Y2=0.0360
r34 24 41 3.59766 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0360 $X2=0.0495 $Y2=0.0360
r35 47 48 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3645
+ $Y=0.0360 $X2=0.3825 $Y2=0.0360
r36 46 47 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0360 $X2=0.3645 $Y2=0.0360
r37 45 46 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.0360 $X2=0.3510 $Y2=0.0360
r38 44 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.0360 $X2=0.3375 $Y2=0.0360
r39 43 44 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3105
+ $Y=0.0360 $X2=0.3240 $Y2=0.0360
r40 42 43 22.0364 $w=1.3e-08 $l=9.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.3105 $Y2=0.0360
r41 40 41 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0675
+ $Y=0.0360 $X2=0.0495 $Y2=0.0360
r42 39 40 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0360 $X2=0.0675 $Y2=0.0360
r43 38 42 22.0364 $w=1.3e-08 $l=9.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1215
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r44 37 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.1215 $Y2=0.0360
r45 22 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.0360 $X2=0.1080 $Y2=0.0360
r46 22 39 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.0360 $X2=0.0810 $Y2=0.0360
r47 14 2 0.958606 $w=2.2e-08 $l=2.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1100 $Y=0.0945 $X2=0.1100 $Y2=0.0725
r48 2 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0540
+ $X2=0.1080 $Y2=0.0360
r49 32 2 0.705882 $w=1.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0980 $Y=0.0725 $X2=0.1100 $Y2=0.0725
r50 17 32 0.264706 $w=1.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0725 $X2=0.0980 $Y2=0.0725
r51 17 2 0.471383 $w=3.35517e-08 $l=3.06472e-08 $layer=N_src_drn
+ $thickness=1e-09 $X=0.0935 $Y=0.0725 $X2=0.1080 $Y2=0.0455
r52 31 29 0.0675676 $w=3.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0455 $X2=0.1225 $Y2=0.0455
r53 2 29 0.391892 $w=3.7e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0455 $X2=0.1225 $Y2=0.0455
r54 2 32 0.441971 $w=3.41429e-08 $l=2.87924e-08 $layer=N_src_drn
+ $thickness=1e-09 $X=0.1080 $Y=0.0455 $X2=0.0980 $Y2=0.0725
r55 13 2 0.391892 $w=3.7e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0455 $X2=0.1080 $Y2=0.0455
r56 30 13 0.0675676 $w=3.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0455 $X2=0.0935 $Y2=0.0455
r57 1 19 1e-05
r58 2 14 1e-05
.ends


*
.SUBCKT AOI21x1_ASAP7_75t_R VSS VDD B A1 A2 Y
*
* VSS VSS
* VDD VDD
* B B
* A1 A1
* A2 A2
* Y Y
*
*

MM4 N_MM4_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3@2 N_MM3@2_d N_MM3@2_g N_MM3@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2@2 N_MM2@2_d N_MM2@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM1@2_g N_MM3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@2 N_MM4@2_d N_MM0@2_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM0 N_MM0_d N_MM4_g N_MM0_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM3@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM2@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@2 N_MM5@2_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1@2 N_MM1@2_d N_MM1@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@2 N_MM0@2_d N_MM0@2_g N_MM0@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AOI21x1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AOI21x1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AOI21x1_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_AOI21x1_ASAP7_75t_R%noxref_12
cc_1 N_noxref_12_1 N_MM0@2_g 0.00344037f
cc_2 N_noxref_12_1 N_Y_16 0.00162515f
x_PM_AOI21x1_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_AOI21x1_ASAP7_75t_R%noxref_10
cc_3 N_noxref_10_1 N_MM4_g 0.00347691f
cc_4 N_noxref_10_1 N_Y_14 0.00159543f
x_PM_AOI21x1_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_AOI21x1_ASAP7_75t_R%noxref_11
cc_5 N_noxref_11_1 N_MM4_g 0.00159475f
cc_6 N_noxref_11_1 N_Y_1 0.000507614f
cc_7 N_noxref_11_1 N_Y_19 0.0374194f
cc_8 N_noxref_11_1 N_noxref_10_1 0.00188935f
x_PM_AOI21x1_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_AOI21x1_ASAP7_75t_R%noxref_13
cc_9 N_noxref_13_1 N_MM0@2_g 0.00158223f
cc_10 N_noxref_13_1 N_Y_4 0.000504597f
cc_11 N_noxref_13_1 N_Y_20 0.0374855f
cc_12 N_noxref_13_1 N_noxref_12_1 0.00189349f
x_PM_AOI21x1_ASAP7_75t_R%NET29__2 VSS N_MM3@2_s N_MM2@2_d N_NET29__2_1
+ PM_AOI21x1_ASAP7_75t_R%NET29__2
cc_13 N_NET29__2_1 N_MM3@2_g 0.0173264f
cc_14 N_NET29__2_1 N_MM2@2_g 0.0173466f
x_PM_AOI21x1_ASAP7_75t_R%A2 VSS A2 N_MM2@2_g N_MM2_g N_A2_1 N_A2_6
+ PM_AOI21x1_ASAP7_75t_R%A2
cc_15 N_A2 N_B_8 0.00595804f
cc_16 N_A2 N_A1_7 0.00139515f
cc_17 N_A2_1 N_A1_1 0.00208878f
cc_18 N_A2_6 N_A1_9 0.00215358f
cc_19 N_MM2@2_g N_MM3@2_g 0.00506534f
cc_20 N_MM2_g N_MM1@2_g 0.00506812f
cc_21 N_A2 N_A1_8 0.00765841f
x_PM_AOI21x1_ASAP7_75t_R%NET29 VSS N_MM2_d N_MM3_s N_NET29_1
+ PM_AOI21x1_ASAP7_75t_R%NET29
cc_22 N_NET29_1 N_MM1@2_g 0.0172733f
cc_23 N_NET29_1 N_MM2_g 0.0173941f
x_PM_AOI21x1_ASAP7_75t_R%NET18 VSS N_MM1@2_d N_MM0@2_s N_MM0_s N_MM1_d N_MM5_d
+ N_MM5@2_d N_NET18_10 N_NET18_1 N_NET18_2 N_NET18_12 N_NET18_3 N_NET18_13
+ N_NET18_11 PM_AOI21x1_ASAP7_75t_R%NET18
cc_24 N_NET18_10 N_MM0@2_g 0.00037116f
cc_25 N_NET18_10 N_B_11 0.000378132f
cc_26 N_NET18_10 N_B_10 0.000396527f
cc_27 N_NET18_10 N_B_8 0.000448469f
cc_28 N_NET18_1 N_B_8 0.000509572f
cc_29 N_NET18_10 N_B_1 0.000604881f
cc_30 N_NET18_2 N_B_8 0.00067507f
cc_31 N_NET18_12 N_B_2 0.000675704f
cc_32 N_NET18_1 N_MM4_g 0.00159091f
cc_33 N_NET18_3 N_MM0@2_g 0.00162601f
cc_34 N_NET18_12 N_MM0@2_g 0.032573f
cc_35 N_NET18_13 N_B_8 0.017166f
cc_36 N_NET18_10 N_MM4_g 0.0343482f
cc_37 N_NET18_12 N_A1_1 0.00063004f
cc_38 N_NET18_3 N_MM1@2_g 0.000900557f
cc_39 N_NET18_1 N_MM3@2_g 0.000924565f
cc_40 N_NET18_10 N_MM3@2_g 0.0327186f
cc_41 N_NET18_12 N_MM1@2_g 0.0353163f
cc_42 N_NET18_11 N_A2_1 0.00195013f
cc_43 N_NET18_2 N_MM2@2_g 0.00196788f
cc_44 N_NET18_11 N_MM2_g 0.0181766f
cc_45 N_NET18_11 N_MM2@2_g 0.049313f
x_PM_AOI21x1_ASAP7_75t_R%B VSS B N_MM4_g N_MM0@2_g N_B_2 N_B_1 N_B_8 N_B_9
+ N_B_7 N_B_11 N_B_10 PM_AOI21x1_ASAP7_75t_R%B
x_PM_AOI21x1_ASAP7_75t_R%A1 VSS A1 N_MM3@2_g N_MM1@2_g N_A1_7 N_A1_2 N_A1_1
+ N_A1_9 N_A1_8 N_A1_10 N_A1_11 PM_AOI21x1_ASAP7_75t_R%A1
cc_46 N_A1_7 N_B_2 0.000935825f
cc_47 N_A1_2 N_B_2 0.00095894f
cc_48 N_A1_1 N_B_1 0.000960942f
cc_49 N_A1_9 N_B_8 0.00243222f
cc_50 N_MM1@2_g N_MM0@2_g 0.00327652f
cc_51 N_MM3@2_g N_MM4_g 0.00328514f
cc_52 N_A1_9 N_B_9 0.00352851f
cc_53 N_A1_7 N_B_7 0.00607897f
x_PM_AOI21x1_ASAP7_75t_R%Y VSS Y N_MM4_d N_MM3@2_d N_MM3_d N_MM4@2_d N_MM0_d
+ N_MM0@2_d N_Y_1 N_Y_4 N_Y_14 N_Y_16 N_Y_19 N_Y_2 N_Y_3 N_Y_22 N_Y_26 N_Y_25
+ N_Y_20 N_Y_23 N_Y_21 N_Y_15 N_Y_13 PM_AOI21x1_ASAP7_75t_R%Y
cc_54 N_Y_1 N_MM0@2_g 0.000230968f
cc_55 N_Y_4 N_MM0@2_g 0.00172255f
cc_56 N_Y_14 N_MM0@2_g 0.000262084f
cc_57 N_Y_16 N_MM0@2_g 0.00556306f
cc_58 N_Y_19 N_MM4_g 0.0537536f
cc_59 N_Y_2 N_B_8 0.000625968f
cc_60 N_Y_2 N_B_1 0.000844484f
cc_61 N_Y_3 N_B_2 0.000913315f
cc_62 N_Y_3 N_MM0@2_g 0.00105828f
cc_63 N_Y_2 N_MM4_g 0.00129831f
cc_64 N_Y_22 N_B_7 0.00137058f
cc_65 N_Y_1 N_MM4_g 0.00147559f
cc_66 N_Y_26 N_B_11 0.00151141f
cc_67 N_Y_25 N_B_10 0.00154315f
cc_68 N_Y_20 N_B_2 0.00178279f
cc_69 N_Y_19 N_B_1 0.00179894f
cc_70 N_Y_23 N_B_9 0.00481891f
cc_71 N_Y_14 N_MM4_g 0.00532681f
cc_72 N_Y_21 N_B_7 0.00735524f
cc_73 N_Y_15 N_MM0@2_g 0.010275f
cc_74 N_Y_13 N_MM4_g 0.0102779f
cc_75 N_Y_20 N_MM0@2_g 0.0546129f
cc_76 N_Y_16 N_MM3@2_g 0.000183843f
cc_77 N_Y_15 N_MM3@2_g 0.00019055f
cc_78 N_Y_2 N_MM3@2_g 0.00217851f
cc_79 N_Y_3 N_MM3@2_g 0.000567495f
cc_80 N_Y_23 N_MM3@2_g 0.000254274f
cc_81 N_Y_2 N_A1_7 0.000683012f
cc_82 N_Y_13 N_A1_1 0.000798329f
cc_83 N_Y_3 N_A1_9 0.000856364f
cc_84 N_Y_15 N_A1_2 0.000913305f
cc_85 N_Y_22 N_A1_10 0.00113933f
cc_86 N_Y_3 N_MM1@2_g 0.00171869f
cc_87 N_Y_22 N_A1_11 0.00189808f
cc_88 N_Y_13 N_MM3@2_g 0.00990963f
cc_89 N_Y_15 N_MM1@2_g 0.00991578f
cc_90 N_Y_22 N_A1_8 0.0128705f
cc_91 N_Y_16 N_MM1@2_g 0.0242707f
cc_92 N_Y_14 N_MM3@2_g 0.0250962f
cc_93 N_Y_26 N_NET18_3 0.000245057f
cc_94 N_Y_19 N_NET18_3 0.00114532f
cc_95 N_Y_20 N_NET18_3 0.00114135f
cc_96 N_Y_1 N_NET18_1 0.00311661f
cc_97 N_Y_25 N_NET18_13 0.000933247f
cc_98 N_Y_4 N_NET18_3 0.00381627f
*END of AOI21x1_ASAP7_75t_R.pxi
.ENDS
** Design:	AOI21xp33_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AOI21xp33_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AOI21xp33_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AOI21xp33_ASAP7_75t_R%noxref_9 VSS 1
c1 1 VSS 0.0319055f
.ends

.subckt PM_AOI21xp33_ASAP7_75t_R%NET29 VSS 2 3 1
c1 1 VSS 0.000853033f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0540 $X2=0.1080 $Y2=0.0540
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0540 $X2=0.1080 $Y2=0.0540
.ends

.subckt PM_AOI21xp33_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.00501026f
.ends

.subckt PM_AOI21xp33_ASAP7_75t_R%A2 VSS 16 3 6 1 9 5
c1 1 VSS 0.00196014f
c2 3 VSS 0.060815f
c3 4 VSS 0.0062534f
c4 5 VSS 0.00279808f
c5 6 VSS 0.0020671f
c6 7 VSS 0.00843887f
c7 8 VSS 0.00127982f
c8 9 VSS 0.00259747f
r1 7 19 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0360 $X2=0.0270 $Y2=0.0540
r2 5 17 5.72052 $w=1.36604e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1660 $X2=0.0270 $Y2=0.1395
r3 5 9 6.28176 $w=1.44063e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1660 $X2=0.0270 $Y2=0.1980
r4 18 19 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0720 $X2=0.0270 $Y2=0.0540
r5 4 8 5.6404 $w=1.39259e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1030 $X2=0.0270 $Y2=0.1300
r6 4 18 7.22888 $w=1.3e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1030 $X2=0.0270 $Y2=0.0720
r7 16 17 0.408178 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1355 $X2=0.0270 $Y2=0.1395
r8 16 8 0.561244 $w=1.8e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1355 $X2=0.0270 $Y2=0.1300
r9 16 15 2.26632 $w=7.16216e-09 $l=1.85607e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1355 $X2=0.0455 $Y2=0.1340
r10 6 13 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.0635
+ $Y=0.1340 $X2=0.0810 $Y2=0.1340
r11 6 15 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0635
+ $Y=0.1340 $X2=0.0455 $Y2=0.1340
r12 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r13 1 13 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1340
.ends

.subckt PM_AOI21xp33_ASAP7_75t_R%B VSS 8 3 1 4
c1 1 VSS 0.00486571f
c2 3 VSS 0.0338359f
c3 4 VSS 0.00368161f
r1 8 4 7.22888 $w=1.3e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1340 $X2=0.1890 $Y2=0.1030
r2 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1340
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AOI21xp33_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.0316694f
.ends

.subckt PM_AOI21xp33_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.00464854f
.ends

.subckt PM_AOI21xp33_ASAP7_75t_R%NET18 VSS 11 21 22 1 9 7 2 8
c1 1 VSS 0.007483f
c2 2 VSS 0.00639586f
c3 7 VSS 0.00323976f
c4 8 VSS 0.00302444f
c5 9 VSS 0.0130636f
r1 22 20 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2160 $X2=0.1765 $Y2=0.2160
r2 2 20 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2160 $X2=0.1765 $Y2=0.2160
r3 8 2 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1620 $Y2=0.2160
r4 21 8 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r5 2 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r6 17 18 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r7 16 17 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.1255
+ $Y=0.2340 $X2=0.1485 $Y2=0.2340
r8 15 16 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1010
+ $Y=0.2340 $X2=0.1255 $Y2=0.2340
r9 14 15 5.13017 $w=1.3e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0790
+ $Y=0.2340 $X2=0.1010 $Y2=0.2340
r10 13 14 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0590
+ $Y=0.2340 $X2=0.0790 $Y2=0.2340
r11 12 13 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0500
+ $Y=0.2340 $X2=0.0590 $Y2=0.2340
r12 9 12 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.2340 $X2=0.0500 $Y2=0.2340
r13 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0500 $Y2=0.2340
r14 11 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r15 7 10 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r16 1 7 1e-05
.ends

.subckt PM_AOI21xp33_ASAP7_75t_R%A1 VSS 4 3 1 5 6
c1 1 VSS 0.00334375f
c2 3 VSS 0.0340695f
c3 4 VSS 0.00229847f
c4 5 VSS 0.00223094f
c5 6 VSS 0.00230359f
r1 6 11 6.28176 $w=1.44063e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1980 $X2=0.1350 $Y2=0.1660
r2 5 10 6.04857 $w=1.44516e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.0720 $X2=0.1350 $Y2=0.1030
r3 4 10 7.22888 $w=1.3e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1340 $X2=0.1350 $Y2=0.1030
r4 4 11 7.46207 $w=1.3e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1340 $X2=0.1350 $Y2=0.1660
r5 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r6 4 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1340
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AOI21xp33_ASAP7_75t_R%Y VSS 25 15 16 33 1 9 7 10 2 8 11
c1 1 VSS 0.00723437f
c2 2 VSS 0.00518232f
c3 7 VSS 0.00391797f
c4 8 VSS 0.00247347f
c5 9 VSS 0.0137504f
c6 10 VSS 0.00491603f
c7 11 VSS 0.0053744f
c8 12 VSS 0.00352772f
r1 8 2 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2160 $X2=0.2140 $Y2=0.2160
r2 33 8 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2160 $X2=0.2015 $Y2=0.2160
r3 2 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2160
+ $X2=0.2160 $Y2=0.2340
r4 30 31 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2295 $Y2=0.2340
r5 11 28 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2430 $Y2=0.2160
r6 11 31 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.2340 $X2=0.2295 $Y2=0.2340
r7 27 28 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2035 $X2=0.2430 $Y2=0.2160
r8 26 27 11.1348 $w=1.3e-08 $l=4.78e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1557 $X2=0.2430 $Y2=0.2035
r9 25 26 10.4352 $w=1.3e-08 $l=4.47e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1110 $X2=0.2430 $Y2=0.1557
r10 25 24 4.83869 $w=1.3e-08 $l=2.08e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1110 $X2=0.2430 $Y2=0.0902
r11 23 24 5.53826 $w=1.3e-08 $l=2.37e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0665 $X2=0.2430 $Y2=0.0902
r12 10 12 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0540 $X2=0.2430 $Y2=0.0360
r13 10 23 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0540 $X2=0.2430 $Y2=0.0665
r14 12 22 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2180 $Y2=0.0360
r15 21 22 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2000
+ $Y=0.0360 $X2=0.2180 $Y2=0.0360
r16 20 21 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.2000 $Y2=0.0360
r17 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1755
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r18 17 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r19 9 17 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r20 1 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r21 16 14 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0540 $X2=0.1765 $Y2=0.0540
r22 1 14 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.0540 $X2=0.1765 $Y2=0.0540
r23 7 1 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1620 $Y2=0.0540
r24 15 7 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
.ends


*
.SUBCKT AOI21xp33_ASAP7_75t_R VSS VDD A2 A1 B Y
*
* VSS VSS
* VDD VDD
* A2 A2
* A1 A1
* B B
* Y Y
*
*

MM2 N_MM2_d N_MM2_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g N_MM3_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM4 N_MM4_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1 N_MM1_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM0 N_MM0_d N_MM4_g N_MM0_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2


*include "AOI21xp33_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AOI21xp33_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AOI21xp33_ASAP7_75t_R%noxref_9 VSS N_noxref_9_1
+ PM_AOI21xp33_ASAP7_75t_R%noxref_9
cc_1 N_noxref_9_1 N_MM2_g 0.00461274f
x_PM_AOI21xp33_ASAP7_75t_R%NET29 VSS N_MM2_d N_MM3_s N_NET29_1
+ PM_AOI21xp33_ASAP7_75t_R%NET29
cc_2 N_NET29_1 N_MM2_g 0.0125189f
cc_3 N_NET29_1 N_MM3_g 0.0125612f
x_PM_AOI21xp33_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_AOI21xp33_ASAP7_75t_R%noxref_10
cc_4 N_noxref_10_1 N_MM2_g 0.00453421f
cc_5 N_noxref_10_1 N_NET18_7 0.0269476f
cc_6 N_noxref_10_1 N_noxref_9_1 0.00204779f
x_PM_AOI21xp33_ASAP7_75t_R%A2 VSS A2 N_MM2_g N_A2_6 N_A2_1 N_A2_9 N_A2_5
+ PM_AOI21xp33_ASAP7_75t_R%A2
x_PM_AOI21xp33_ASAP7_75t_R%B VSS B N_MM4_g N_B_1 N_B_4
+ PM_AOI21xp33_ASAP7_75t_R%B
cc_7 N_B_1 N_A1_1 0.00263773f
cc_8 N_B_4 N_A1 0.00452621f
cc_9 N_MM4_g N_MM3_g 0.00810841f
x_PM_AOI21xp33_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_AOI21xp33_ASAP7_75t_R%noxref_11
cc_10 N_noxref_11_1 N_MM4_g 0.00367842f
cc_11 N_noxref_11_1 N_Y_7 0.00117334f
x_PM_AOI21xp33_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_AOI21xp33_ASAP7_75t_R%noxref_12
cc_12 N_noxref_12_1 N_MM4_g 0.00367842f
cc_13 N_noxref_12_1 N_Y_8 0.0282032f
cc_14 N_noxref_12_1 N_noxref_11_1 0.00205576f
x_PM_AOI21xp33_ASAP7_75t_R%NET18 VSS N_MM5_d N_MM1_d N_MM0_s N_NET18_1
+ N_NET18_9 N_NET18_7 N_NET18_2 N_NET18_8 PM_AOI21xp33_ASAP7_75t_R%NET18
cc_15 N_NET18_1 N_A2_9 0.000385761f
cc_16 N_NET18_1 N_A2_5 0.000401184f
cc_17 N_NET18_1 N_MM2_g 0.00115648f
cc_18 N_NET18_9 N_A2_9 0.00340531f
cc_19 N_NET18_7 N_MM2_g 0.0255973f
cc_20 N_NET18_2 N_MM3_g 0.000709987f
cc_21 N_NET18_9 N_A1_6 0.00414715f
cc_22 N_NET18_8 N_MM3_g 0.0256156f
cc_23 N_NET18_2 N_MM4_g 0.000700762f
cc_24 N_NET18_2 N_B_4 0.000775329f
cc_25 N_NET18_8 N_MM4_g 0.0253613f
x_PM_AOI21xp33_ASAP7_75t_R%A1 VSS A1 N_MM3_g N_A1_1 N_A1_5 N_A1_6
+ PM_AOI21xp33_ASAP7_75t_R%A1
cc_26 N_A1_1 N_A2_6 0.000481014f
cc_27 N_A1_5 N_A2_6 0.000645773f
cc_28 N_A1_1 N_A2_1 0.00253491f
cc_29 N_A1 N_A2_6 0.00276317f
cc_30 N_MM3_g N_MM2_g 0.0101401f
x_PM_AOI21xp33_ASAP7_75t_R%Y VSS Y N_MM3_d N_MM4_d N_MM0_d N_Y_1 N_Y_9 N_Y_7
+ N_Y_10 N_Y_2 N_Y_8 N_Y_11 PM_AOI21xp33_ASAP7_75t_R%Y
cc_31 N_Y_1 N_A1 0.000605656f
cc_32 N_Y_1 N_MM3_g 0.000975355f
cc_33 N_Y_9 N_A1_5 0.00412534f
cc_34 N_Y_7 N_MM3_g 0.0265844f
cc_35 N_Y_10 N_B_1 0.000588369f
cc_36 N_Y_1 N_MM4_g 0.000726967f
cc_37 N_Y_2 N_MM4_g 0.000748702f
cc_38 N_Y_8 N_B_1 0.00074952f
cc_39 N_Y_9 N_B_4 0.00107108f
cc_40 N_Y_8 N_MM4_g 0.0108853f
cc_41 N_Y_10 N_B_4 0.0079171f
cc_42 N_Y_7 N_MM4_g 0.0399554f
cc_43 N_Y_2 N_NET18_8 0.00042317f
cc_44 N_Y_11 N_NET18_9 0.000932493f
cc_45 N_Y_2 N_NET18_2 0.00313894f
*END of AOI21xp33_ASAP7_75t_R.pxi
.ENDS
** Design:	AOI21xp5_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AOI21xp5_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AOI21xp5_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AOI21xp5_ASAP7_75t_R%NET29 VSS 2 3 1
c1 1 VSS 0.00103056f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_AOI21xp5_ASAP7_75t_R%noxref_9 VSS 1
c1 1 VSS 0.0419366f
.ends

.subckt PM_AOI21xp5_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.00644175f
.ends

.subckt PM_AOI21xp5_ASAP7_75t_R%A2 VSS 14 3 1 6 5
c1 1 VSS 0.00483435f
c2 3 VSS 0.0822377f
c3 4 VSS 0.011865f
c4 5 VSS 0.00525235f
c5 6 VSS 0.0030299f
c6 7 VSS 0.00168591f
r1 5 15 7.00306 $w=1.35469e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1715 $X2=0.0270 $Y2=0.1395
r2 4 7 6.92294 $w=1.37692e-08 $l=3.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0975 $X2=0.0270 $Y2=0.1300
r3 14 15 0.408178 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1355 $X2=0.0270 $Y2=0.1395
r4 14 7 0.561244 $w=1.8e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1355 $X2=0.0270 $Y2=0.1300
r5 14 13 0.517402 $w=3.18182e-09 $l=1.11018e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1355 $X2=0.0380 $Y2=0.1340
r6 6 11 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.0560
+ $Y=0.1340 $X2=0.0810 $Y2=0.1340
r7 6 13 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0560
+ $Y=0.1340 $X2=0.0380 $Y2=0.1340
r8 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r9 1 11 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1340
.ends

.subckt PM_AOI21xp5_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.00479001f
.ends

.subckt PM_AOI21xp5_ASAP7_75t_R%A1 VSS 4 3 1
c1 1 VSS 0.00715394f
c2 3 VSS 0.0459573f
c3 4 VSS 0.00540515f
r1 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r2 4 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1340
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AOI21xp5_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.0316168f
.ends

.subckt PM_AOI21xp5_ASAP7_75t_R%B VSS 8 3 4 1
c1 1 VSS 0.00656732f
c2 3 VSS 0.0346058f
c3 4 VSS 0.00465988f
r1 8 4 8.51143 $w=1.3e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1340 $X2=0.1890 $Y2=0.0975
r2 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1340
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AOI21xp5_ASAP7_75t_R%NET18 VSS 11 19 22 7 9 1 2 8
c1 1 VSS 0.00798563f
c2 2 VSS 0.00719456f
c3 7 VSS 0.0036853f
c4 8 VSS 0.00327837f
c5 9 VSS 0.0130172f
r1 22 21 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r2 20 21 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1720 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r3 2 20 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1600 $Y=0.2025 $X2=0.1720 $Y2=0.2025
r4 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1600 $Y2=0.2025
r5 19 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r6 2 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r7 16 17 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r8 15 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1485 $Y2=0.2340
r9 14 15 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1105
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r10 13 14 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0790
+ $Y=0.2340 $X2=0.1105 $Y2=0.2340
r11 12 13 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2340 $X2=0.0790 $Y2=0.2340
r12 9 12 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r13 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r14 11 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r15 7 10 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r16 1 7 1e-05
.ends

.subckt PM_AOI21xp5_ASAP7_75t_R%Y VSS 31 17 18 38 8 11 1 7 2 10 12 13
c1 1 VSS 0.00858257f
c2 2 VSS 0.00527033f
c3 7 VSS 0.00327942f
c4 8 VSS 0.000579196f
c5 9 VSS 6.55989e-20
c6 10 VSS 0.00237883f
c7 11 VSS 0.0100671f
c8 12 VSS 0.00429692f
c9 13 VSS 0.0058853f
c10 14 VSS 0.0034103f
r1 10 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2140 $Y2=0.2025
r2 38 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r3 2 35 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.2340
r4 35 36 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2295 $Y2=0.2340
r5 13 33 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.2340 $X2=0.2430 $Y2=0.2125
r6 13 36 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.2340 $X2=0.2295 $Y2=0.2340
r7 32 33 13.2335 $w=1.3e-08 $l=5.68e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1557 $X2=0.2430 $Y2=0.2125
r8 31 32 10.4352 $w=1.3e-08 $l=4.47e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1110 $X2=0.2430 $Y2=0.1557
r9 31 30 4.83869 $w=1.3e-08 $l=2.08e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1110 $X2=0.2430 $Y2=0.0902
r10 12 14 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0575 $X2=0.2430 $Y2=0.0360
r11 12 30 7.63696 $w=1.3e-08 $l=3.27e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0575 $X2=0.2430 $Y2=0.0902
r12 14 29 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2180 $Y2=0.0360
r13 28 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2000
+ $Y=0.0360 $X2=0.2180 $Y2=0.0360
r14 27 28 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.2000 $Y2=0.0360
r15 26 27 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1755
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r16 24 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r17 11 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r18 8 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0945 $X2=0.1600 $Y2=0.0945
r19 1 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r20 20 21 0.264706 $w=1.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1720 $Y=0.0725 $X2=0.1765 $Y2=0.0725
r21 1 20 0.705882 $w=1.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1600 $Y=0.0725 $X2=0.1720 $Y2=0.0725
r22 9 1 0.735294 $w=1.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0725 $X2=0.1600 $Y2=0.0725
r23 18 16 0.0675676 $w=3.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0455 $X2=0.1765 $Y2=0.0455
r24 1 16 0.391892 $w=3.7e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.0455 $X2=0.1765 $Y2=0.0455
r25 1 21 0.471383 $w=3.35517e-08 $l=3.06472e-08 $layer=N_src_drn
+ $thickness=1e-09 $X=0.1620 $Y=0.0455 $X2=0.1765 $Y2=0.0725
r26 7 1 0.391892 $w=3.7e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0455 $X2=0.1620 $Y2=0.0455
r27 17 7 0.0675676 $w=3.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0455 $X2=0.1475 $Y2=0.0455
.ends


*
.SUBCKT AOI21xp5_ASAP7_75t_R VSS VDD A2 A1 B Y
*
* VSS VSS
* VDD VDD
* A2 A2
* A1 A1
* B B
* Y Y
*
*

MM2 N_MM2_d N_MM2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g N_MM3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM4_g N_MM0_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AOI21xp5_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AOI21xp5_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AOI21xp5_ASAP7_75t_R%NET29 VSS N_MM2_d N_MM3_s N_NET29_1
+ PM_AOI21xp5_ASAP7_75t_R%NET29
cc_1 N_NET29_1 N_MM2_g 0.0174231f
cc_2 N_NET29_1 N_MM3_g 0.0172649f
x_PM_AOI21xp5_ASAP7_75t_R%noxref_9 VSS N_noxref_9_1
+ PM_AOI21xp5_ASAP7_75t_R%noxref_9
cc_3 N_noxref_9_1 N_MM2_g 0.00217537f
cc_4 N_noxref_9_1 N_NET18_7 0.000481873f
x_PM_AOI21xp5_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_AOI21xp5_ASAP7_75t_R%noxref_10
cc_5 N_noxref_10_1 N_MM2_g 0.00208607f
cc_6 N_noxref_10_1 N_NET18_7 0.0361025f
cc_7 N_noxref_10_1 N_noxref_9_1 0.00176185f
x_PM_AOI21xp5_ASAP7_75t_R%A2 VSS A2 N_MM2_g N_A2_1 N_A2_6 N_A2_5
+ PM_AOI21xp5_ASAP7_75t_R%A2
x_PM_AOI21xp5_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_AOI21xp5_ASAP7_75t_R%noxref_12
cc_8 N_noxref_12_1 N_MM4_g 0.00159491f
cc_9 N_noxref_12_1 N_Y_10 0.0381663f
cc_10 N_noxref_12_1 N_noxref_11_1 0.00188743f
x_PM_AOI21xp5_ASAP7_75t_R%A1 VSS A1 N_MM3_g N_A1_1 PM_AOI21xp5_ASAP7_75t_R%A1
cc_11 N_A1_1 N_A2_1 0.00122691f
cc_12 N_A1 N_A2_6 0.00287678f
cc_13 N_MM3_g N_MM2_g 0.00641531f
x_PM_AOI21xp5_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_AOI21xp5_ASAP7_75t_R%noxref_11
cc_14 N_noxref_11_1 N_MM4_g 0.0034589f
cc_15 N_noxref_11_1 N_Y_8 0.0016031f
x_PM_AOI21xp5_ASAP7_75t_R%B VSS B N_MM4_g N_B_4 N_B_1 PM_AOI21xp5_ASAP7_75t_R%B
cc_16 N_MM4_g N_MM3_g 0.00328019f
cc_17 N_B_4 N_A1 0.00629039f
x_PM_AOI21xp5_ASAP7_75t_R%NET18 VSS N_MM5_d N_MM1_d N_MM0_s N_NET18_7 N_NET18_9
+ N_NET18_1 N_NET18_2 N_NET18_8 PM_AOI21xp5_ASAP7_75t_R%NET18
cc_18 N_NET18_7 N_A2_1 0.00080399f
cc_19 N_NET18_9 N_A2_5 0.00096699f
cc_20 N_NET18_1 N_A2_5 0.00149875f
cc_21 N_NET18_1 N_MM2_g 0.00182775f
cc_22 N_NET18_7 N_MM2_g 0.0350386f
cc_23 N_NET18_2 N_MM3_g 0.00114917f
cc_24 N_NET18_9 N_A1 0.00116222f
cc_25 N_NET18_2 N_A1 0.0017867f
cc_26 N_NET18_8 N_MM3_g 0.0346724f
cc_27 N_NET18_8 N_B_1 0.0007348f
cc_28 N_NET18_2 N_B_4 0.00095414f
cc_29 N_NET18_2 N_MM4_g 0.00119135f
cc_30 N_NET18_8 N_MM4_g 0.034156f
x_PM_AOI21xp5_ASAP7_75t_R%Y VSS Y N_MM3_d N_MM4_d N_MM0_d N_Y_8 N_Y_11 N_Y_1
+ N_Y_7 N_Y_2 N_Y_10 N_Y_12 N_Y_13 PM_AOI21xp5_ASAP7_75t_R%Y
cc_31 N_Y_8 N_A1_1 0.000639132f
cc_32 N_Y_11 N_A1 0.000713349f
cc_33 N_Y_1 N_MM3_g 0.00157565f
cc_34 N_Y_1 N_A1 0.00158332f
cc_35 N_Y_7 N_MM3_g 0.00994985f
cc_36 N_Y_8 N_MM3_g 0.0255929f
cc_37 N_Y_1 N_B_1 0.000818091f
cc_38 N_Y_11 N_B_4 0.00107165f
cc_39 N_Y_1 N_MM4_g 0.00132487f
cc_40 N_Y_2 N_MM4_g 0.00138975f
cc_41 N_Y_10 N_B_1 0.00163784f
cc_42 N_Y_8 N_MM4_g 0.00531385f
cc_43 N_Y_12 N_B_4 0.00777949f
cc_44 N_Y_7 N_MM4_g 0.0103293f
cc_45 N_Y_10 N_MM4_g 0.0553628f
cc_46 N_Y_10 N_NET18_8 0.000595311f
cc_47 N_Y_13 N_NET18_9 0.000818844f
cc_48 N_Y_2 N_NET18_2 0.00418874f
*END of AOI21xp5_ASAP7_75t_R.pxi
.ENDS
** Design:	AOI221x1_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AOI221x1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AOI221x1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AOI221x1_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00698823f
.ends

.subckt PM_AOI221x1_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.0422353f
.ends

.subckt PM_AOI221x1_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.00653999f
.ends

.subckt PM_AOI221x1_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.04247f
.ends

.subckt PM_AOI221x1_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.00568398f
.ends

.subckt PM_AOI221x1_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.0051558f
.ends

.subckt PM_AOI221x1_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.00581542f
.ends

.subckt PM_AOI221x1_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.00512619f
.ends

.subckt PM_AOI221x1_ASAP7_75t_R%NET16 VSS 19 22 36 39 41 43 1 13 2 14 3 15 4 16
+ 17
c1 1 VSS 0.00459699f
c2 2 VSS 0.00441473f
c3 3 VSS 0.00494538f
c4 4 VSS 0.00542406f
c5 13 VSS 0.00222699f
c6 14 VSS 0.00221208f
c7 15 VSS 0.00227035f
c8 16 VSS 0.00231389f
c9 17 VSS 0.0338634f
r1 16 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.2025 $X2=0.7000 $Y2=0.2025
r2 43 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.2025 $X2=0.6875 $Y2=0.2025
r3 41 40 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.2025 $X2=0.6085 $Y2=0.2025
r4 15 40 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5960 $Y=0.2025 $X2=0.6085 $Y2=0.2025
r5 39 38 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r6 2 38 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4340 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r7 35 2 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4220 $Y=0.2025 $X2=0.4340 $Y2=0.2025
r8 14 35 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4220 $Y2=0.2025
r9 36 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r10 4 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7020 $Y=0.2025
+ $X2=0.7020 $Y2=0.2340
r11 3 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2025
+ $X2=0.5940 $Y2=0.2340
r12 2 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.2340
r13 32 33 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.6635
+ $Y=0.2340 $X2=0.7020 $Y2=0.2340
r14 31 32 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.6185
+ $Y=0.2340 $X2=0.6635 $Y2=0.2340
r15 30 31 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.2340 $X2=0.6185 $Y2=0.2340
r16 29 30 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5805
+ $Y=0.2340 $X2=0.5940 $Y2=0.2340
r17 28 29 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5575
+ $Y=0.2340 $X2=0.5805 $Y2=0.2340
r18 27 28 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5195
+ $Y=0.2340 $X2=0.5575 $Y2=0.2340
r19 26 27 11.4263 $w=1.3e-08 $l=4.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4705
+ $Y=0.2340 $X2=0.5195 $Y2=0.2340
r20 25 26 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4705 $Y2=0.2340
r21 24 25 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.4320 $Y2=0.2340
r22 23 24 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r23 17 23 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3125
+ $Y=0.2340 $X2=0.3240 $Y2=0.2340
r24 1 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.2340
r25 22 21 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r26 20 21 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3340 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r27 1 20 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3220 $Y=0.2025 $X2=0.3340 $Y2=0.2025
r28 13 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3220 $Y2=0.2025
r29 19 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r30 3 15 1e-05
.ends

.subckt PM_AOI221x1_ASAP7_75t_R%C VSS 26 3 4 6 1 9 7 8
c1 1 VSS 0.00646441f
c2 3 VSS 0.0344462f
c3 4 VSS 0.0354695f
c4 5 VSS 0.00274882f
c5 6 VSS 0.00307973f
c6 7 VSS 0.00310064f
c7 8 VSS 0.00407208f
c8 9 VSS 0.00475586f
c9 10 VSS 0.00260513f
r1 28 29 0.280622 $w=1.8e-08 $l=2.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.5710
+ $Y=0.1980 $X2=0.5737 $Y2=0.1980
r2 9 28 0.6888 $w=1.8e-08 $l=6.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.5642
+ $Y=0.1980 $X2=0.5710 $Y2=0.1980
r3 26 9 0.754373 $w=1.76296e-08 $l=9.90404e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.1885 $X2=0.5642 $Y2=0.1980
r4 26 29 0.346195 $w=1.70909e-08 $l=1.1625e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.1885 $X2=0.5737 $Y2=0.1980
r5 26 25 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1885 $X2=0.5670 $Y2=0.1795
r6 24 25 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1620 $X2=0.5670 $Y2=0.1795
r7 6 10 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.1485 $X2=0.5670 $Y2=0.1350
r8 6 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1485 $X2=0.5670 $Y2=0.1620
r9 5 10 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1125 $X2=0.5670 $Y2=0.1350
r10 5 8 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1125 $X2=0.5670 $Y2=0.0900
r11 4 19 2.92627 $w=1.245e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.6750
+ $Y=0.1350 $X2=0.6750 $Y2=0.1345
r12 7 21 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.1350 $X2=0.6210 $Y2=0.1350
r13 7 10 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5940 $Y=0.1350 $X2=0.5670 $Y2=0.1350
r14 17 19 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6625 $Y=0.1345 $X2=0.6750 $Y2=0.1345
r15 16 17 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6480 $Y=0.1345 $X2=0.6625 $Y2=0.1345
r16 15 16 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6335 $Y=0.1345 $X2=0.6480 $Y2=0.1345
r17 13 15 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.6305 $Y=0.1345 $X2=0.6335 $Y2=0.1345
r18 12 13 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.6210
+ $Y=0.1345 $X2=0.6305 $Y2=0.1345
r19 12 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6210 $Y=0.1345
+ $X2=0.6210 $Y2=0.1350
r20 1 12 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.6115
+ $Y=0.1345 $X2=0.6210 $Y2=0.1345
r21 1 14 0.721303 $w=1.75333e-08 $l=1.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.6115 $Y=0.1345 $X2=0.6100 $Y2=0.1345
r22 3 12 2.66511 $w=1.29895e-07 $l=5e-10 $layer=LIG $thickness=5.22105e-08
+ $X=0.6210 $Y=0.1350 $X2=0.6210 $Y2=0.1345
r23 3 14 0.905388 $w=2.07755e-07 $l=1.10114e-08 $layer=LIG
+ $thickness=5.52727e-08 $X=0.6210 $Y=0.1350 $X2=0.6100 $Y2=0.1345
r24 3 15 1.79147 $w=1.8466e-07 $l=1.251e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.6210 $Y=0.1350 $X2=0.6335 $Y2=0.1345
.ends

.subckt PM_AOI221x1_ASAP7_75t_R%A1 VSS 21 3 4 1 5 7
c1 1 VSS 0.011128f
c2 3 VSS 0.0463416f
c3 4 VSS 0.0456562f
c4 5 VSS 0.00485802f
c5 6 VSS 0.00872662f
c6 7 VSS 0.00410901f
r1 7 24 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1620 $X2=0.1890 $Y2=0.1485
r2 6 22 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.1890 $Y2=0.0540
r3 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1485
r4 21 20 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0807 $X2=0.1890 $Y2=0.0717
r5 20 22 4.13912 $w=1.3e-08 $l=1.77e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0717 $X2=0.1890 $Y2=0.0540
r6 18 19 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0812 $X2=0.1890 $Y2=0.0902
r7 21 18 0.116595 $w=1.3e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0807 $X2=0.1890 $Y2=0.0812
r8 5 19 5.18847 $w=1.3e-08 $l=2.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1125 $X2=0.1890 $Y2=0.0902
r9 5 23 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1125 $X2=0.1890 $Y2=0.1350
r10 3 14 2.66511 $w=1.29895e-07 $l=5e-10 $layer=LIG $thickness=5.22105e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1890 $Y2=0.1345
r11 14 15 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1890
+ $Y=0.1345 $X2=0.1985 $Y2=0.1345
r12 14 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1345
+ $X2=0.1890 $Y2=0.1350
r13 11 15 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.2015 $Y=0.1345 $X2=0.1985 $Y2=0.1345
r14 10 11 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2160 $Y=0.1345 $X2=0.2015 $Y2=0.1345
r15 9 10 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2305 $Y=0.1345 $X2=0.2160 $Y2=0.1345
r16 4 1 2.92627 $w=1.245e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1345
r17 1 9 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2430 $Y=0.1345 $X2=0.2305 $Y2=0.1345
r18 1 17 3.05464 $w=2.15326e-08 $l=1.07e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2430 $Y=0.1345 $X2=0.2537 $Y2=0.1345
r19 4 9 1.79147 $w=1.8466e-07 $l=1.251e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2305 $Y2=0.1345
r20 4 17 0.757708 $w=2.1223e-07 $l=1.07117e-08 $layer=LIG
+ $thickness=5.54419e-08 $X=0.2430 $Y=0.1350 $X2=0.2537 $Y2=0.1345
.ends

.subckt PM_AOI221x1_ASAP7_75t_R%NET10 VSS 24 25 54 55 58 59 61 63 16 2 1 21 17
+ 18 3 19 4 20 5
c1 1 VSS 0.00738517f
c2 2 VSS 0.00852577f
c3 3 VSS 0.00604919f
c4 4 VSS 0.0028608f
c5 5 VSS 0.00448335f
c6 16 VSS 0.00371737f
c7 17 VSS 0.0044414f
c8 18 VSS 0.00339895f
c9 19 VSS 0.0021759f
c10 20 VSS 0.00288182f
c11 21 VSS 0.0141173f
r1 20 5 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4840 $Y2=0.2025
r2 63 20 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r3 61 60 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r4 16 60 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r5 59 57 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r6 2 57 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r7 17 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r8 58 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r9 55 53 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r10 3 53 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r11 18 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r12 54 18 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r13 5 49 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2025
+ $X2=0.4820 $Y2=0.1980
r14 1 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0580 $Y2=0.1980
r15 2 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1660 $Y2=0.1980
r16 3 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2740 $Y2=0.1980
r17 48 49 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4725
+ $Y=0.1980 $X2=0.4820 $Y2=0.1980
r18 47 48 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1980 $X2=0.4725 $Y2=0.1980
r19 46 47 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4205
+ $Y=0.1980 $X2=0.4590 $Y2=0.1980
r20 42 43 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0580
+ $Y=0.1980 $X2=0.0675 $Y2=0.1980
r21 41 43 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1980 $X2=0.0675 $Y2=0.1980
r22 40 41 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1195
+ $Y=0.1980 $X2=0.0810 $Y2=0.1980
r23 38 39 1.39914 $w=1.3e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.1510
+ $Y=0.1980 $X2=0.1570 $Y2=0.1980
r24 38 40 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1510
+ $Y=0.1980 $X2=0.1195 $Y2=0.1980
r25 36 37 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1660
+ $Y=0.1980 $X2=0.1755 $Y2=0.1980
r26 36 39 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1660
+ $Y=0.1980 $X2=0.1570 $Y2=0.1980
r27 35 37 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.1985
+ $Y=0.1980 $X2=0.1755 $Y2=0.1980
r28 34 35 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2365
+ $Y=0.1980 $X2=0.1985 $Y2=0.1980
r29 32 33 1.51573 $w=1.3e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2585
+ $Y=0.1980 $X2=0.2650 $Y2=0.1980
r30 32 34 5.13018 $w=1.3e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2585
+ $Y=0.1980 $X2=0.2365 $Y2=0.1980
r31 30 31 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2740
+ $Y=0.1980 $X2=0.2925 $Y2=0.1980
r32 30 33 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2740
+ $Y=0.1980 $X2=0.2650 $Y2=0.1980
r33 29 31 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3080
+ $Y=0.1980 $X2=0.2925 $Y2=0.1980
r34 28 29 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3175
+ $Y=0.1980 $X2=0.3080 $Y2=0.1980
r35 27 46 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3890
+ $Y=0.1980 $X2=0.4205 $Y2=0.1980
r36 26 27 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.1980 $X2=0.3890 $Y2=0.1980
r37 21 26 7.22888 $w=1.3e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3470
+ $Y=0.1980 $X2=0.3780 $Y2=0.1980
r38 21 28 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.3470
+ $Y=0.1980 $X2=0.3175 $Y2=0.1980
r39 4 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.1980
r40 25 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r41 4 23 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r42 19 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3780 $Y2=0.2025
r43 24 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r44 1 16 1e-05
.ends

.subckt PM_AOI221x1_ASAP7_75t_R%NET24 VSS 11 19 8 2 1 3 9 5
c1 1 VSS 0.00624962f
c2 2 VSS 0.00279319f
c3 3 VSS 0.000330353f
c4 5 VSS 0.00313315f
c5 8 VSS 0.00333916f
c6 9 VSS 0.00216875f
r1 19 18 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r2 9 18 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2180 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r3 3 5 16.8928 $w=2.18031e-08 $l=3.2e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.2160 $Y=0.0895 $X2=0.2160 $Y2=0.0575
r4 5 16 12.2208 $w=2.36037e-08 $l=2.53e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.2160 $Y=0.0575 $X2=0.1907 $Y2=0.0575
r5 15 16 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.1757 $Y=0.0575 $X2=0.1907 $Y2=0.0575
r6 14 15 6.46718 $w=2.32e-08 $l=1.37e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.1620 $Y=0.0575 $X2=0.1757 $Y2=0.0575
r7 13 14 6.46718 $w=2.32e-08 $l=1.38e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.1482 $Y=0.0575 $X2=0.1620 $Y2=0.0575
r8 2 1 12.2208 $w=2.36037e-08 $l=2.52e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.1332 $Y=0.0575 $X2=0.1080 $Y2=0.0575
r9 2 13 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.1332
+ $Y=0.0575 $X2=0.1482 $Y2=0.0575
r10 8 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0675 $X2=0.1060 $Y2=0.0675
r11 11 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.0935 $Y2=0.0675
r12 3 9 1e-05
r13 5 9 1e-05
.ends

.subckt PM_AOI221x1_ASAP7_75t_R%A2 VSS 20 3 4 6 8 9 1
c1 1 VSS 0.0106982f
c2 3 VSS 0.0825507f
c3 4 VSS 0.0451753f
c4 5 VSS 0.00524902f
c5 6 VSS 0.00334706f
c6 7 VSS 0.00883761f
c7 8 VSS 0.00276679f
c8 9 VSS 0.00304719f
r1 8 25 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0625 $Y=0.1620 $X2=0.0810 $Y2=0.1620
r2 5 9 10.3626 $w=1.39091e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0855 $X2=0.0810 $Y2=0.1350
r3 5 7 10.3626 $w=1.39091e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0855 $X2=0.0810 $Y2=0.0360
r4 24 25 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1485 $X2=0.0810 $Y2=0.1620
r5 9 24 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0810 $Y2=0.1485
r6 21 22 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1150
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r7 20 21 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1035
+ $Y=0.1350 $X2=0.1150 $Y2=0.1350
r8 20 6 1.63233 $w=1.3e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1035
+ $Y=0.1350 $X2=0.0965 $Y2=0.1350
r9 6 9 2.43413 $w=1.59032e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0965 $Y=0.1350 $X2=0.0810 $Y2=0.1350
r10 4 17 2.66511 $w=1.29895e-07 $l=5e-10 $layer=LIG $thickness=5.22105e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1350 $Y2=0.1345
r11 17 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1345
+ $X2=0.1350 $Y2=0.1350
r12 16 17 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1255
+ $Y=0.1345 $X2=0.1350 $Y2=0.1345
r13 14 16 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1345 $X2=0.1255 $Y2=0.1345
r14 13 14 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1345 $X2=0.1225 $Y2=0.1345
r15 12 13 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1345 $X2=0.1080 $Y2=0.1345
r16 3 1 2.92627 $w=1.245e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1345
r17 1 11 3.05464 $w=2.15326e-08 $l=1.08e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0810 $Y=0.1345 $X2=0.0702 $Y2=0.1345
r18 1 12 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0810 $Y=0.1345 $X2=0.0935 $Y2=0.1345
r19 3 11 0.757708 $w=2.1223e-07 $l=1.08116e-08 $layer=LIG
+ $thickness=5.54419e-08 $X=0.0810 $Y=0.1350 $X2=0.0702 $Y2=0.1345
r20 3 12 1.79147 $w=1.8466e-07 $l=1.251e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1345
.ends

.subckt PM_AOI221x1_ASAP7_75t_R%NET23 VSS 11 17 4 2 8 5 9 3 1
c1 1 VSS 0.00324906f
c2 2 VSS 0.00074038f
c3 3 VSS 0.00497979f
c4 4 VSS 0.000136357f
c5 5 VSS 0.00114041f
c6 8 VSS 0.00226837f
c7 9 VSS 0.00346552f
r1 17 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r2 9 16 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4340 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r3 3 5 21.3436 $w=2.22923e-08 $l=4.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4320 $Y=0.0540 $X2=0.4320 $Y2=0.0945
r4 5 15 10.5221 $w=2.51178e-08 $l=2.53e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.4320 $Y=0.0945 $X2=0.4067 $Y2=0.0945
r5 14 15 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.3917 $Y=0.0945 $X2=0.4067 $Y2=0.0945
r6 13 14 6.46718 $w=2.32e-08 $l=1.37e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.3780 $Y=0.0945 $X2=0.3917 $Y2=0.0945
r7 12 13 6.46718 $w=2.32e-08 $l=1.38e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.3642 $Y=0.0945 $X2=0.3780 $Y2=0.0945
r8 2 4 10.5221 $w=2.51178e-08 $l=2.52e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.3492 $Y=0.0945 $X2=0.3240 $Y2=0.0945
r9 2 12 7.05511 $w=2.32e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08 $X=0.3492
+ $Y=0.0945 $X2=0.3642 $Y2=0.0945
r10 1 4 21.3436 $w=2.22923e-08 $l=4.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.3240 $Y=0.0540 $X2=0.3240 $Y2=0.0945
r11 8 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3220 $Y2=0.0675
r12 11 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r13 3 9 1e-05
r14 5 9 1e-05
r15 1 4 1e-05
.ends

.subckt PM_AOI221x1_ASAP7_75t_R%Y VSS 42 20 21 38 50 53 13 1 10 14 2 11 3 15 12
+ 17
c1 1 VSS 0.00435626f
c2 2 VSS 0.0063744f
c3 3 VSS 0.00289474f
c4 10 VSS 0.00225522f
c5 11 VSS 0.00321104f
c6 12 VSS 0.00225408f
c7 13 VSS 0.0272786f
c8 14 VSS 0.000796135f
c9 15 VSS 0.00227928f
c10 16 VSS 0.00193772f
c11 17 VSS 0.000800369f
r1 53 52 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.2025 $X2=0.6625 $Y2=0.2025
r2 51 52 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6580 $Y=0.2025 $X2=0.6625 $Y2=0.2025
r3 3 51 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6460 $Y=0.2025 $X2=0.6580 $Y2=0.2025
r4 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.2025 $X2=0.6460 $Y2=0.2025
r5 50 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.2025 $X2=0.6335 $Y2=0.2025
r6 3 46 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.2025
+ $X2=0.6480 $Y2=0.1980
r7 46 47 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.6480
+ $Y=0.1980 $X2=0.6865 $Y2=0.1980
r8 14 17 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7180 $Y=0.1980 $X2=0.7290 $Y2=0.1980
r9 14 47 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.7180
+ $Y=0.1980 $X2=0.6865 $Y2=0.1980
r10 17 44 5.69636 $w=1.58e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1980 $X2=0.7290 $Y2=0.1665
r11 43 44 6.41272 $w=1.3e-08 $l=2.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1390 $X2=0.7290 $Y2=0.1665
r12 42 43 1.28254 $w=1.3e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1335 $X2=0.7290 $Y2=0.1390
r13 42 41 0.932759 $w=1.3e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1335 $X2=0.7290 $Y2=0.1295
r14 40 41 3.96423 $w=1.3e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1125 $X2=0.7290 $Y2=0.1295
r15 39 40 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.0900 $X2=0.7290 $Y2=0.1125
r16 15 16 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.0720 $X2=0.7290 $Y2=0.0540
r17 15 39 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.0720 $X2=0.7290 $Y2=0.0900
r18 38 37 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.0540 $X2=0.6085 $Y2=0.0540
r19 11 37 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5960 $Y=0.0540 $X2=0.6085 $Y2=0.0540
r20 16 36 10.2436 $w=1.38824e-08 $l=5.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.0540 $X2=0.6780 $Y2=0.0540
r21 2 34 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0540
+ $X2=0.5940 $Y2=0.0540
r22 35 36 13.6416 $w=1.3e-08 $l=5.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.6195
+ $Y=0.0540 $X2=0.6780 $Y2=0.0540
r23 34 35 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0540 $X2=0.6195 $Y2=0.0540
r24 33 34 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5805
+ $Y=0.0540 $X2=0.5940 $Y2=0.0540
r25 32 33 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5575
+ $Y=0.0540 $X2=0.5805 $Y2=0.0540
r26 31 32 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5195
+ $Y=0.0540 $X2=0.5575 $Y2=0.0540
r27 30 31 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.4935
+ $Y=0.0540 $X2=0.5195 $Y2=0.0540
r28 29 30 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.4775
+ $Y=0.0540 $X2=0.4935 $Y2=0.0540
r29 28 29 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4495
+ $Y=0.0540 $X2=0.4775 $Y2=0.0540
r30 27 28 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4110
+ $Y=0.0540 $X2=0.4495 $Y2=0.0540
r31 26 27 12.3591 $w=1.3e-08 $l=5.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.3580
+ $Y=0.0540 $X2=0.4110 $Y2=0.0540
r32 25 26 12.0093 $w=1.3e-08 $l=5.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3065
+ $Y=0.0540 $X2=0.3580 $Y2=0.0540
r33 24 25 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.2835
+ $Y=0.0540 $X2=0.3065 $Y2=0.0540
r34 23 24 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2740
+ $Y=0.0540 $X2=0.2835 $Y2=0.0540
r35 22 23 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2650
+ $Y=0.0540 $X2=0.2740 $Y2=0.0540
r36 13 22 1.51573 $w=1.3e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2585
+ $Y=0.0540 $X2=0.2650 $Y2=0.0540
r37 1 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2740 $Y2=0.0540
r38 21 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r39 1 19 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r40 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r41 20 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
r42 2 11 1e-05
.ends

.subckt PM_AOI221x1_ASAP7_75t_R%B2 VSS 24 3 4 9 8 1 5 7
c1 1 VSS 0.0079322f
c2 3 VSS 0.00809255f
c3 4 VSS 0.0458475f
c4 5 VSS 0.00363788f
c5 6 VSS 0.00366804f
c6 7 VSS 0.00427642f
c7 8 VSS 0.00349737f
c8 9 VSS 0.00440134f
r1 9 25 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4775 $Y=0.1620 $X2=0.4590 $Y2=0.1620
r2 6 8 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1125 $X2=0.4590 $Y2=0.1350
r3 6 7 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1125 $X2=0.4590 $Y2=0.0900
r4 24 25 1.03499 $w=1.77368e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1525 $X2=0.4590 $Y2=0.1620
r5 24 23 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1525 $X2=0.4590 $Y2=0.1480
r6 8 21 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4405 $Y2=0.1350
r7 8 23 1.85116 $w=1.64615e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4590 $Y2=0.1480
r8 4 17 2.92627 $w=1.245e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1345
r9 20 21 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4225
+ $Y=0.1350 $X2=0.4405 $Y2=0.1350
r10 19 20 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4225 $Y2=0.1350
r11 5 19 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3935
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r12 15 17 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4465 $Y=0.1345 $X2=0.4590 $Y2=0.1345
r13 14 15 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4320 $Y=0.1345 $X2=0.4465 $Y2=0.1345
r14 13 14 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4175 $Y=0.1345 $X2=0.4320 $Y2=0.1345
r15 11 13 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.4145 $Y=0.1345 $X2=0.4175 $Y2=0.1345
r16 10 11 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.4050
+ $Y=0.1345 $X2=0.4145 $Y2=0.1345
r17 10 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1345
+ $X2=0.4050 $Y2=0.1350
r18 1 10 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.3955
+ $Y=0.1345 $X2=0.4050 $Y2=0.1345
r19 1 12 0.573622 $w=1.798e-08 $l=1.3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.3955 $Y=0.1345 $X2=0.3942 $Y2=0.1345
r20 3 10 2.66511 $w=1.29895e-07 $l=5e-10 $layer=LIG $thickness=5.22105e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4050 $Y2=0.1345
r21 3 12 0.757708 $w=2.1223e-07 $l=1.08116e-08 $layer=LIG
+ $thickness=5.54419e-08 $X=0.4050 $Y=0.1350 $X2=0.3942 $Y2=0.1345
r22 3 13 1.79147 $w=1.8466e-07 $l=1.251e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4175 $Y2=0.1345
.ends

.subckt PM_AOI221x1_ASAP7_75t_R%B1 VSS 18 3 4 1 6 7
c1 1 VSS 0.00859562f
c2 3 VSS 0.00874289f
c3 4 VSS 0.00932962f
c4 5 VSS 0.00467625f
c5 6 VSS 0.0047238f
c6 7 VSS 0.00463315f
r1 6 21 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1620 $X2=0.2970 $Y2=0.1485
r2 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1485
r3 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1215 $X2=0.2970 $Y2=0.1350
r4 18 19 1.16595 $w=1.3e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1165 $X2=0.2970 $Y2=0.1215
r5 18 5 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1165 $X2=0.2970 $Y2=0.1075
r6 5 7 2.90051 $w=1.55714e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1075 $X2=0.2970 $Y2=0.0900
r7 3 13 2.66511 $w=1.29895e-07 $l=5e-10 $layer=LIG $thickness=5.22105e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2970 $Y2=0.1345
r8 13 14 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2970
+ $Y=0.1345 $X2=0.3065 $Y2=0.1345
r9 13 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1345
+ $X2=0.2970 $Y2=0.1350
r10 10 14 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.3095 $Y=0.1345 $X2=0.3065 $Y2=0.1345
r11 9 10 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3240 $Y=0.1345 $X2=0.3095 $Y2=0.1345
r12 8 9 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08 $X=0.3385
+ $Y=0.1345 $X2=0.3240 $Y2=0.1345
r13 4 1 2.92627 $w=1.245e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1345
r14 1 8 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3510 $Y=0.1345 $X2=0.3385 $Y2=0.1345
r15 1 16 3.05464 $w=2.15326e-08 $l=1.07e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3510 $Y=0.1345 $X2=0.3617 $Y2=0.1345
r16 4 8 1.79147 $w=1.8466e-07 $l=1.251e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.3510 $Y=0.1350 $X2=0.3385 $Y2=0.1345
r17 4 16 0.757708 $w=2.1223e-07 $l=1.07117e-08 $layer=LIG
+ $thickness=5.54419e-08 $X=0.3510 $Y=0.1350 $X2=0.3617 $Y2=0.1345
.ends


*
.SUBCKT AOI221x1_ASAP7_75t_R VSS VDD A2 A1 B1 B2 C Y
*
* VSS VSS
* VDD VDD
* A2 A2
* A1 A1
* B1 B1
* B2 B2
* C C
* Y Y
*
*

MM0 N_MM0_d N_MM0_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM26 N_MM26_d N_MM26_g N_MM26_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM27 N_MM27_d N_MM32@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM28 N_MM28_d N_MM1_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM31 N_MM31_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM31@2 N_MM31@2_d N_MM31@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM29 N_MM29_d N_MM29_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM29@2 N_MM29@2_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM30 N_MM30_d N_MM26_g N_MM30_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM30@2 N_MM30@2_d N_MM30@2_g N_MM30@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM32 N_MM32_d N_MM32_g N_MM32_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM32@2 N_MM32@2_d N_MM32@2_g N_MM32@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1@2 N_MM1@2_d N_MM1@2_g N_MM1@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AOI221x1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AOI221x1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AOI221x1_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_AOI221x1_ASAP7_75t_R%noxref_14
cc_1 N_noxref_14_1 N_MM0_g 0.00165724f
cc_2 N_noxref_14_1 N_NET10_16 0.035967f
cc_3 N_noxref_14_1 N_noxref_13_1 0.00178885f
x_PM_AOI221x1_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_AOI221x1_ASAP7_75t_R%noxref_13
cc_4 N_noxref_13_1 N_MM0_g 0.00174663f
cc_5 N_noxref_13_1 N_NET10_16 0.000582407f
x_PM_AOI221x1_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_AOI221x1_ASAP7_75t_R%noxref_16
cc_6 N_noxref_16_1 N_MM32@2_g 0.00141107f
cc_7 N_noxref_16_1 N_NET10_20 0.0354243f
cc_8 N_noxref_16_1 N_NET16_14 0.000680919f
cc_9 N_noxref_16_1 N_noxref_15_1 0.0012324f
x_PM_AOI221x1_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_AOI221x1_ASAP7_75t_R%noxref_15
cc_10 N_noxref_15_1 N_MM32@2_g 0.00142358f
cc_11 N_noxref_15_1 N_Y_11 0.000566579f
x_PM_AOI221x1_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_AOI221x1_ASAP7_75t_R%noxref_20
cc_12 N_noxref_20_1 N_MM1@2_g 0.00164244f
cc_13 N_noxref_20_1 N_NET16_16 0.0363769f
cc_14 N_noxref_20_1 N_Y_12 0.000794815f
cc_15 N_noxref_20_1 N_noxref_19_1 0.00194363f
x_PM_AOI221x1_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_AOI221x1_ASAP7_75t_R%noxref_19
cc_16 N_noxref_19_1 N_MM1@2_g 0.00911342f
cc_17 N_noxref_19_1 N_NET16_16 0.000628487f
cc_18 N_noxref_19_1 N_Y_15 0.00137938f
x_PM_AOI221x1_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_AOI221x1_ASAP7_75t_R%noxref_18
cc_19 N_noxref_18_1 N_MM1_g 0.00181329f
cc_20 N_noxref_18_1 N_NET10_20 0.000551683f
cc_21 N_noxref_18_1 N_NET16_15 0.0361931f
cc_22 N_noxref_18_1 N_noxref_16_1 0.00766118f
cc_23 N_noxref_18_1 N_noxref_17_1 0.00135208f
x_PM_AOI221x1_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_AOI221x1_ASAP7_75t_R%noxref_17
cc_24 N_noxref_17_1 N_MM1_g 0.00369609f
cc_25 N_noxref_17_1 N_NET16_15 0.000467881f
cc_26 N_noxref_17_1 N_Y_11 0.0268711f
cc_27 N_noxref_17_1 N_noxref_15_1 0.0076993f
cc_28 N_noxref_17_1 N_noxref_16_1 0.000470588f
x_PM_AOI221x1_ASAP7_75t_R%NET16 VSS N_MM30_d N_MM30@2_d N_MM32_d N_MM32@2_d
+ N_MM1_s N_MM1@2_s N_NET16_1 N_NET16_13 N_NET16_2 N_NET16_14 N_NET16_3
+ N_NET16_15 N_NET16_4 N_NET16_16 N_NET16_17 PM_AOI221x1_ASAP7_75t_R%NET16
cc_29 N_NET16_1 N_MM30@2_g 0.00192579f
cc_30 N_NET16_13 N_B1_1 0.00197356f
cc_31 N_NET16_13 N_MM26_g 0.0184532f
cc_32 N_NET16_13 N_MM30@2_g 0.0495505f
cc_33 N_NET16_2 N_MM32@2_g 0.00229966f
cc_34 N_NET16_14 N_B2_1 0.00195459f
cc_35 N_NET16_14 N_MM32_g 0.0184514f
cc_36 N_NET16_14 N_MM32@2_g 0.0498282f
cc_37 N_NET16_3 N_MM1@2_g 0.000395567f
cc_38 N_NET16_15 N_MM1@2_g 0.000472433f
cc_39 N_NET16_3 N_C_6 0.000725661f
cc_40 N_NET16_4 N_MM1@2_g 0.000877269f
cc_41 N_NET16_16 N_C_1 0.00175054f
cc_42 N_NET16_3 N_MM1_g 0.00187209f
cc_43 N_NET16_17 N_C_9 0.0050814f
cc_44 N_NET16_15 N_MM1_g 0.0338335f
cc_45 N_NET16_16 N_MM1@2_g 0.0350325f
cc_46 N_NET16_17 N_NET10_5 0.000507381f
cc_47 N_NET16_13 N_NET10_18 0.000554657f
cc_48 N_NET16_17 N_NET10_4 0.000636627f
cc_49 N_NET16_14 N_NET10_20 0.00176701f
cc_50 N_NET16_2 N_NET10_21 0.000742733f
cc_51 N_NET16_1 N_NET10_21 0.000798874f
cc_52 N_NET16_14 N_NET10_19 0.00111597f
cc_53 N_NET16_13 N_NET10_19 0.00112716f
cc_54 N_NET16_1 N_NET10_3 0.00125007f
cc_55 N_NET16_2 N_NET10_4 0.0027651f
cc_56 N_NET16_1 N_NET10_4 0.00309537f
cc_57 N_NET16_2 N_NET10_5 0.00485264f
cc_58 N_NET16_17 N_NET10_21 0.0188155f
x_PM_AOI221x1_ASAP7_75t_R%C VSS C N_MM1_g N_MM1@2_g N_C_6 N_C_1 N_C_9 N_C_7
+ N_C_8 PM_AOI221x1_ASAP7_75t_R%C
x_PM_AOI221x1_ASAP7_75t_R%A1 VSS A1 N_MM29_g N_MM2_g N_A1_1 N_A1_5 N_A1_7
+ PM_AOI221x1_ASAP7_75t_R%A1
cc_59 N_A1_1 N_MM31@2_g 0.00126141f
cc_60 N_A1_5 N_A2_6 0.00219988f
cc_61 N_MM29_g N_MM31@2_g 0.012604f
x_PM_AOI221x1_ASAP7_75t_R%NET10 VSS N_MM30@2_s N_MM32_s N_MM29@2_d N_MM30_s
+ N_MM31@2_d N_MM29_d N_MM31_d N_MM32@2_s N_NET10_16 N_NET10_2 N_NET10_1
+ N_NET10_21 N_NET10_17 N_NET10_18 N_NET10_3 N_NET10_19 N_NET10_4 N_NET10_20
+ N_NET10_5 PM_AOI221x1_ASAP7_75t_R%NET10
cc_62 N_NET10_16 N_MM31@2_g 0.000486044f
cc_63 N_NET10_2 N_MM31@2_g 0.000888256f
cc_64 N_NET10_1 N_MM0_g 0.00117472f
cc_65 N_NET10_21 N_A2_8 0.00122013f
cc_66 N_NET10_21 N_A2_9 0.00152144f
cc_67 N_NET10_17 N_A2_1 0.00166221f
cc_68 N_NET10_21 N_A2_6 0.00374488f
cc_69 N_NET10_16 N_MM0_g 0.0330138f
cc_70 N_NET10_17 N_MM31@2_g 0.0345507f
cc_71 N_NET10_18 N_MM29_g 0.000433916f
cc_72 N_NET10_3 N_MM29_g 0.000748884f
cc_73 N_NET10_2 N_MM29_g 0.000925197f
cc_74 N_NET10_18 N_A1_1 0.00163975f
cc_75 N_NET10_21 N_A1_7 0.00489091f
cc_76 N_NET10_18 N_MM2_g 0.0329087f
cc_77 N_NET10_17 N_MM29_g 0.0345422f
cc_78 N_NET10_21 N_MM26_g 0.000378751f
cc_79 N_NET10_19 N_MM26_g 0.000436529f
cc_80 N_NET10_4 N_MM30@2_g 0.000734818f
cc_81 N_NET10_3 N_MM26_g 0.00101816f
cc_82 N_NET10_19 N_B1_1 0.00169321f
cc_83 N_NET10_21 N_B1_6 0.00501115f
cc_84 N_NET10_19 N_MM30@2_g 0.033028f
cc_85 N_NET10_18 N_MM26_g 0.0342466f
cc_86 N_NET10_20 N_MM32_g 0.000433142f
cc_87 N_NET10_4 N_MM32_g 0.000889514f
cc_88 N_NET10_5 N_MM32@2_g 0.00112113f
cc_89 N_NET10_21 N_B2_9 0.00133733f
cc_90 N_NET10_21 N_B2_8 0.0015622f
cc_91 N_NET10_20 N_B2_1 0.00161123f
cc_92 N_NET10_21 N_B2_5 0.00401735f
cc_93 N_NET10_20 N_MM32@2_g 0.0330693f
cc_94 N_NET10_19 N_MM32_g 0.0344459f
x_PM_AOI221x1_ASAP7_75t_R%NET24 VSS N_MM0_d N_MM2_s N_NET24_8 N_NET24_2
+ N_NET24_1 N_NET24_3 N_NET24_9 N_NET24_5 PM_AOI221x1_ASAP7_75t_R%NET24
cc_95 N_NET24_8 N_MM0_g 0.030108f
cc_96 N_NET24_2 N_MM31@2_g 0.00166199f
cc_97 N_NET24_1 N_MM31@2_g 0.00222637f
cc_98 N_NET24_8 N_A2_1 0.00228645f
cc_99 N_NET24_8 N_MM31@2_g 0.0429116f
cc_100 N_NET24_3 N_MM2_g 0.00208461f
cc_101 N_NET24_9 N_A1_1 0.00230841f
cc_102 N_NET24_2 N_MM29_g 0.0023653f
cc_103 N_NET24_9 N_MM29_g 0.0197658f
cc_104 N_NET24_9 N_MM2_g 0.054134f
cc_105 N_NET24_5 N_Y_10 0.00112127f
cc_106 N_NET24_5 N_Y_1 0.00361376f
x_PM_AOI221x1_ASAP7_75t_R%A2 VSS A2 N_MM0_g N_MM31@2_g N_A2_6 N_A2_8 N_A2_9
+ N_A2_1 PM_AOI221x1_ASAP7_75t_R%A2
x_PM_AOI221x1_ASAP7_75t_R%NET23 VSS N_MM26_s N_MM27_d N_NET23_4 N_NET23_2
+ N_NET23_8 N_NET23_5 N_NET23_9 N_NET23_3 N_NET23_1
+ PM_AOI221x1_ASAP7_75t_R%NET23
cc_107 N_NET23_4 N_B1_1 0.00149361f
cc_108 N_NET23_2 N_B1_1 0.00282223f
cc_109 N_NET23_8 N_B1_1 0.00303965f
cc_110 N_NET23_8 N_MM26_g 0.029635f
cc_111 N_NET23_8 N_MM30@2_g 0.0433244f
cc_112 N_NET23_5 N_B2_1 0.0015712f
cc_113 N_NET23_9 N_B2_1 0.00300215f
cc_114 N_NET23_2 N_B2_1 0.00310159f
cc_115 N_NET23_9 N_MM32_g 0.0198103f
cc_116 N_NET23_9 N_MM32@2_g 0.0536929f
cc_117 N_NET23_3 N_Y_10 0.00114718f
cc_118 N_NET23_3 N_Y_1 0.000698608f
cc_119 N_NET23_1 N_Y_1 0.00278083f
cc_120 N_NET23_3 N_Y_13 0.00429118f
x_PM_AOI221x1_ASAP7_75t_R%Y VSS Y N_MM2_d N_MM26_d N_MM28_d N_MM1_d N_MM1@2_d
+ N_Y_13 N_Y_1 N_Y_10 N_Y_14 N_Y_2 N_Y_11 N_Y_3 N_Y_15 N_Y_12 N_Y_17
+ PM_AOI221x1_ASAP7_75t_R%Y
cc_121 N_Y_13 N_MM2_g 0.000958906f
cc_122 N_Y_1 N_MM2_g 0.000876147f
cc_123 N_Y_10 N_MM2_g 0.0353825f
cc_124 N_Y_1 N_MM26_g 0.00165457f
cc_125 N_Y_13 N_B1_7 0.00219874f
cc_126 N_Y_13 N_B1_1 0.00267578f
cc_127 N_Y_10 N_MM26_g 0.035691f
cc_128 N_Y_13 N_B2_7 0.00666399f
cc_129 N_Y_14 N_MM1_g 0.000277596f
cc_130 N_Y_2 N_MM1_g 0.00119438f
cc_131 N_Y_11 N_MM1_g 0.0112106f
cc_132 N_Y_13 N_MM1_g 0.000437109f
cc_133 N_Y_3 N_C_1 0.000751506f
cc_134 N_Y_15 N_C_1 0.000846244f
cc_135 N_Y_12 N_MM1@2_g 0.0497593f
cc_136 N_Y_3 N_MM1@2_g 0.0018822f
cc_137 N_Y_14 N_C_7 0.00246292f
cc_138 N_Y_12 N_C_1 0.00332993f
cc_139 N_Y_13 N_C_8 0.00665277f
cc_140 N_Y_12 N_MM1_g 0.0328302f
cc_141 N_Y_12 N_NET16_15 0.00059529f
cc_142 N_Y_17 N_NET16_17 0.000619663f
cc_143 N_Y_14 N_NET16_4 0.000683076f
cc_144 N_Y_12 N_NET16_16 0.00182151f
cc_145 N_Y_3 N_NET16_17 0.000789005f
cc_146 N_Y_15 N_NET16_4 0.000815345f
cc_147 N_Y_3 N_NET16_3 0.00141678f
cc_148 N_Y_3 N_NET16_4 0.0053536f
cc_149 N_Y_14 N_NET16_17 0.00925767f
x_PM_AOI221x1_ASAP7_75t_R%B2 VSS B2 N_MM32_g N_MM32@2_g N_B2_9 N_B2_8 N_B2_1
+ N_B2_5 N_B2_7 PM_AOI221x1_ASAP7_75t_R%B2
cc_150 N_MM32_g N_MM30@2_g 0.0122737f
x_PM_AOI221x1_ASAP7_75t_R%B1 VSS B1 N_MM26_g N_MM30@2_g N_B1_1 N_B1_6 N_B1_7
+ PM_AOI221x1_ASAP7_75t_R%B1
cc_151 N_MM26_g N_MM2_g 0.00608829f
*END of AOI221x1_ASAP7_75t_R.pxi
.ENDS
** Design:	AOI221xp5_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AOI221xp5_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AOI221xp5_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AOI221xp5_ASAP7_75t_R%NET23 VSS 2 3 1
c1 1 VSS 0.000848583f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0540 $X2=0.1080 $Y2=0.0540
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0540 $X2=0.1080 $Y2=0.0540
.ends

.subckt PM_AOI221xp5_ASAP7_75t_R%NET24 VSS 2 3 1
c1 1 VSS 0.000855142f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0540 $X2=0.2700 $Y2=0.0540
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0540 $X2=0.2700 $Y2=0.0540
.ends

.subckt PM_AOI221xp5_ASAP7_75t_R%B2 VSS 6 3 1 4
c1 1 VSS 0.00553028f
c2 3 VSS 0.0353397f
c3 4 VSS 0.00422091f
r1 7 8 4.02252 $w=1.3e-08 $l=1.73e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1177 $X2=0.1350 $Y2=0.1350
r2 6 7 2.04041 $w=1.3e-08 $l=8.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1090 $X2=0.1350 $Y2=0.1177
r3 6 4 4.6055 $w=1.3e-08 $l=1.98e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1090 $X2=0.1350 $Y2=0.0892
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AOI221xp5_ASAP7_75t_R%B1 VSS 8 3 1 4
c1 1 VSS 0.00665986f
c2 3 VSS 0.0085276f
c3 4 VSS 0.00423482f
r1 8 7 0.524677 $w=1.3e-08 $l=2.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1480 $X2=0.0810 $Y2=0.1457
r2 6 7 2.50679 $w=1.3e-08 $l=1.07e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1457
r3 4 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0980 $X2=0.0810 $Y2=0.1350
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r5 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AOI221xp5_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00476099f
.ends

.subckt PM_AOI221xp5_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00555622f
.ends

.subckt PM_AOI221xp5_ASAP7_75t_R%Y VSS 35 19 39 40 48 49 2 1 15 14 12 10 13 3
+ 11 17
c1 1 VSS 0.00550983f
c2 2 VSS 0.00282553f
c3 3 VSS 0.00779554f
c4 10 VSS 0.00257204f
c5 11 VSS 0.00371314f
c6 12 VSS 0.0021541f
c7 13 VSS 0.00205115f
c8 14 VSS 0.0189996f
c9 15 VSS 0.000791706f
c10 16 VSS 0.00307376f
c11 17 VSS 0.000770888f
r1 49 47 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r2 2 47 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r3 12 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r4 48 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
r5 2 44 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.1980
r6 43 44 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.1980 $X2=0.1080 $Y2=0.1980
r7 42 43 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1980 $X2=0.0945 $Y2=0.1980
r8 41 42 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.0560
+ $Y=0.1980 $X2=0.0810 $Y2=0.1980
r9 15 17 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0380 $Y=0.1980 $X2=0.0270 $Y2=0.1980
r10 15 41 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0380
+ $Y=0.1980 $X2=0.0560 $Y2=0.1980
r11 17 36 2.37341 $w=1.8113e-08 $l=1.73e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1980 $X2=0.0270 $Y2=0.1807
r12 40 38 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0540 $X2=0.2305 $Y2=0.0540
r13 3 38 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.0540 $X2=0.2305 $Y2=0.0540
r14 11 3 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0540 $X2=0.2160 $Y2=0.0540
r15 39 11 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0540 $X2=0.2015 $Y2=0.0540
r16 35 36 2.04041 $w=1.3e-08 $l=8.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1720 $X2=0.0270 $Y2=0.1807
r17 35 34 0.991056 $w=1.3e-08 $l=4.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1720 $X2=0.0270 $Y2=0.1677
r18 33 34 11.8344 $w=1.3e-08 $l=5.07e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1170 $X2=0.0270 $Y2=0.1677
r19 13 16 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0575 $X2=0.0270 $Y2=0.0360
r20 13 33 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0575 $X2=0.0270 $Y2=0.1170
r21 3 31 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0540
+ $X2=0.2160 $Y2=0.0360
r22 30 31 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2040
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r23 29 30 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1995
+ $Y=0.0360 $X2=0.2040 $Y2=0.0360
r24 28 29 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.1995 $Y2=0.0360
r25 27 28 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1780
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r26 26 27 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1600
+ $Y=0.0360 $X2=0.1780 $Y2=0.0360
r27 25 26 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1600 $Y2=0.0360
r28 24 25 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1245
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r29 23 24 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1065
+ $Y=0.0360 $X2=0.1245 $Y2=0.0360
r30 22 23 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0360 $X2=0.1065 $Y2=0.0360
r31 21 22 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0675
+ $Y=0.0360 $X2=0.0810 $Y2=0.0360
r32 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.0360 $X2=0.0675 $Y2=0.0360
r33 14 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r34 14 16 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0405 $Y=0.0360 $X2=0.0270 $Y2=0.0360
r35 1 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0540 $Y2=0.0360
r36 19 18 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r37 10 18 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r38 1 10 1e-05
.ends

.subckt PM_AOI221xp5_ASAP7_75t_R%NET16 VSS 11 21 22 7 1 8 2 9
c1 1 VSS 0.00520287f
c2 2 VSS 0.00461746f
c3 7 VSS 0.0022178f
c4 8 VSS 0.00213415f
c5 9 VSS 0.0120826f
r1 22 20 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r2 2 20 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r4 21 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r5 2 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r6 16 17 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r7 15 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1485 $Y2=0.2340
r8 14 15 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1245
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r9 13 14 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0930
+ $Y=0.2340 $X2=0.1245 $Y2=0.2340
r10 12 13 9.0944 $w=1.3e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2340 $X2=0.0930 $Y2=0.2340
r11 9 12 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r12 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r13 11 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r14 7 10 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r15 1 7 1e-05
.ends

.subckt PM_AOI221xp5_ASAP7_75t_R%C VSS 6 3 1 4
c1 1 VSS 0.00658235f
c2 3 VSS 0.0347966f
c3 4 VSS 0.00463168f
r1 7 8 2.39019 $w=1.3e-08 $l=1.03e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1247 $X2=0.1890 $Y2=0.1350
r2 6 7 0.408082 $w=1.3e-08 $l=1.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1230 $X2=0.1890 $Y2=0.1247
r3 6 4 6.23783 $w=1.3e-08 $l=2.68e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1230 $X2=0.1890 $Y2=0.0962
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AOI221xp5_ASAP7_75t_R%A1 VSS 6 3 1 4
c1 1 VSS 0.00676546f
c2 3 VSS 0.0457645f
c3 4 VSS 0.0041058f
r1 7 8 6.23783 $w=1.3e-08 $l=2.68e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1082 $X2=0.2430 $Y2=0.1350
r2 6 7 4.25571 $w=1.3e-08 $l=1.82e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0900 $X2=0.2430 $Y2=0.1082
r3 6 4 2.39019 $w=1.3e-08 $l=1.03e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0900 $X2=0.2430 $Y2=0.0797
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AOI221xp5_ASAP7_75t_R%A2 VSS 6 3 1 4
c1 1 VSS 0.00361444f
c2 3 VSS 0.0714007f
c3 4 VSS 0.0149724f
r1 7 8 2.39019 $w=1.3e-08 $l=1.03e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1247 $X2=0.2970 $Y2=0.1350
r2 6 7 0.408082 $w=1.3e-08 $l=1.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1230 $X2=0.2970 $Y2=0.1247
r3 6 4 6.23783 $w=1.3e-08 $l=2.68e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1230 $X2=0.2970 $Y2=0.0962
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_AOI221xp5_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.00638752f
.ends

.subckt PM_AOI221xp5_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.032019f
.ends

.subckt PM_AOI221xp5_ASAP7_75t_R%NET012 VSS 12 13 24 7 1 9 8 2
c1 1 VSS 0.0061757f
c2 2 VSS 0.00720264f
c3 7 VSS 0.00336125f
c4 8 VSS 0.00353499f
c5 9 VSS 0.0066394f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3220 $Y2=0.2025
r2 24 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r3 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3230 $Y2=0.1980
r4 20 21 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.3100
+ $Y=0.1980 $X2=0.3230 $Y2=0.1980
r5 19 20 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1980 $X2=0.3100 $Y2=0.1980
r6 18 19 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1980 $X2=0.2970 $Y2=0.1980
r7 17 18 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1980 $X2=0.2700 $Y2=0.1980
r8 16 17 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2320
+ $Y=0.1980 $X2=0.2430 $Y2=0.1980
r9 15 16 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2275
+ $Y=0.1980 $X2=0.2320 $Y2=0.1980
r10 14 15 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1980 $X2=0.2275 $Y2=0.1980
r11 9 14 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2040
+ $Y=0.1980 $X2=0.2160 $Y2=0.1980
r12 1 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.1980
r13 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r14 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r15 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r16 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
.ends


*
.SUBCKT AOI221xp5_ASAP7_75t_R VSS VDD B1 B2 C A1 A2 Y
*
* VSS VSS
* VDD VDD
* B1 B1
* B2 B2
* C C
* A1 A1
* A2 A2
* Y Y
*
*

MM26 N_MM26_d N_MM26_g N_MM26_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM27 N_MM27_d N_MM27_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM28 N_MM28_d N_MM28_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2 N_MM2_d N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM0 N_MM0_d N_MM0_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM30 N_MM30_d N_MM26_g N_MM30_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM32 N_MM32_d N_MM27_g N_MM32_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM28_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM29 N_MM29_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM31 N_MM31_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AOI221xp5_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AOI221xp5_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AOI221xp5_ASAP7_75t_R%NET23 VSS N_MM26_s N_MM27_d N_NET23_1
+ PM_AOI221xp5_ASAP7_75t_R%NET23
cc_1 N_NET23_1 N_MM26_g 0.0125009f
cc_2 N_NET23_1 N_MM27_g 0.0125359f
x_PM_AOI221xp5_ASAP7_75t_R%NET24 VSS N_MM2_s N_MM0_d N_NET24_1
+ PM_AOI221xp5_ASAP7_75t_R%NET24
cc_3 N_NET24_1 N_MM2_g 0.0125064f
cc_4 N_NET24_1 N_MM0_g 0.0125668f
x_PM_AOI221xp5_ASAP7_75t_R%B2 VSS B2 N_MM27_g N_B2_1 N_B2_4
+ PM_AOI221xp5_ASAP7_75t_R%B2
cc_5 N_B2_1 N_B1_1 0.00134947f
cc_6 N_B2_4 N_B1_4 0.00336995f
cc_7 N_MM27_g N_MM26_g 0.0075452f
x_PM_AOI221xp5_ASAP7_75t_R%B1 VSS B1 N_MM26_g N_B1_1 N_B1_4
+ PM_AOI221xp5_ASAP7_75t_R%B1
x_PM_AOI221xp5_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_AOI221xp5_ASAP7_75t_R%noxref_13
cc_8 N_noxref_13_1 N_MM26_g 0.00350437f
cc_9 N_noxref_13_1 N_Y_10 0.0279048f
cc_10 N_noxref_13_1 N_NET16_7 0.000582539f
x_PM_AOI221xp5_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_AOI221xp5_ASAP7_75t_R%noxref_14
cc_11 N_noxref_14_1 N_MM26_g 0.00159641f
cc_12 N_noxref_14_1 N_Y_12 0.000865415f
cc_13 N_noxref_14_1 N_NET16_7 0.0364547f
cc_14 N_noxref_14_1 N_noxref_13_1 0.0018973f
x_PM_AOI221xp5_ASAP7_75t_R%Y VSS Y N_MM26_d N_MM28_d N_MM2_d N_MM30_s N_MM32_s
+ N_Y_2 N_Y_1 N_Y_15 N_Y_14 N_Y_12 N_Y_10 N_Y_13 N_Y_3 N_Y_11 N_Y_17
+ PM_AOI221xp5_ASAP7_75t_R%Y
cc_15 N_Y_2 N_B1_1 0.000761567f
cc_16 N_Y_2 N_MM26_g 0.000899131f
cc_17 N_Y_1 N_MM26_g 0.000934162f
cc_18 N_Y_15 N_B1_4 0.00112495f
cc_19 N_Y_14 N_B1_4 0.00117558f
cc_20 N_Y_12 N_B1_1 0.00132331f
cc_21 N_Y_10 N_MM26_g 0.0107945f
cc_22 N_Y_13 N_B1_4 0.00652699f
cc_23 N_Y_12 N_MM26_g 0.0490817f
cc_24 N_Y_15 N_B2_4 0.00057505f
cc_25 N_Y_12 N_B2_1 0.000736981f
cc_26 N_Y_2 N_MM27_g 0.000916383f
cc_27 N_Y_14 N_B2_4 0.00131176f
cc_28 N_Y_2 N_B2_4 0.00218789f
cc_29 N_Y_12 N_MM27_g 0.0357115f
cc_30 N_Y_14 N_C_4 0.00112274f
cc_31 N_Y_3 N_C_4 0.00157406f
cc_32 N_Y_11 N_MM28_g 0.0258972f
cc_33 N_Y_3 N_MM2_g 0.000931816f
cc_34 N_Y_3 N_A1_4 0.00110923f
cc_35 N_Y_11 N_MM2_g 0.0262695f
x_PM_AOI221xp5_ASAP7_75t_R%NET16 VSS N_MM30_d N_MM32_d N_MM1_s N_NET16_7
+ N_NET16_1 N_NET16_8 N_NET16_2 N_NET16_9 PM_AOI221xp5_ASAP7_75t_R%NET16
cc_36 N_NET16_7 N_B1_1 0.000856925f
cc_37 N_NET16_1 N_MM26_g 0.00103933f
cc_38 N_NET16_7 N_MM26_g 0.0346023f
cc_39 N_NET16_8 N_B2_1 0.000603535f
cc_40 N_NET16_2 N_MM27_g 0.000976859f
cc_41 N_NET16_8 N_MM27_g 0.0347317f
cc_42 N_NET16_8 N_C_1 0.000682219f
cc_43 N_NET16_2 N_MM28_g 0.000977192f
cc_44 N_NET16_8 N_MM28_g 0.0345613f
cc_45 N_NET16_8 N_Y_15 0.000564963f
cc_46 N_NET16_9 N_Y_17 0.000623936f
cc_47 N_NET16_1 N_Y_13 0.000704809f
cc_48 N_NET16_7 N_Y_12 0.000713147f
cc_49 N_NET16_9 N_Y_2 0.000797009f
cc_50 N_NET16_8 N_Y_12 0.00112624f
cc_51 N_NET16_1 N_Y_2 0.00241506f
cc_52 N_NET16_2 N_Y_2 0.00420877f
cc_53 N_NET16_9 N_Y_15 0.00963944f
x_PM_AOI221xp5_ASAP7_75t_R%C VSS C N_MM28_g N_C_1 N_C_4
+ PM_AOI221xp5_ASAP7_75t_R%C
cc_54 N_C_1 N_B2_1 0.00126825f
cc_55 N_C_4 N_B2_4 0.0033729f
cc_56 N_MM28_g N_MM27_g 0.0063088f
x_PM_AOI221xp5_ASAP7_75t_R%A1 VSS A1 N_MM2_g N_A1_1 N_A1_4
+ PM_AOI221xp5_ASAP7_75t_R%A1
cc_57 N_A1_1 N_C_1 0.00117857f
cc_58 N_A1_4 N_C_4 0.00340132f
cc_59 N_MM2_g N_MM28_g 0.00622566f
x_PM_AOI221xp5_ASAP7_75t_R%A2 VSS A2 N_MM0_g N_A2_1 N_A2_4
+ PM_AOI221xp5_ASAP7_75t_R%A2
cc_60 N_A2_1 N_A1_1 0.00131213f
cc_61 N_A2_4 N_A1_4 0.00404958f
cc_62 N_MM0_g N_MM2_g 0.00771124f
x_PM_AOI221xp5_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_AOI221xp5_ASAP7_75t_R%noxref_16
cc_63 N_noxref_16_1 N_MM0_g 0.00174125f
cc_64 N_noxref_16_1 N_NET012_8 0.0362603f
cc_65 N_noxref_16_1 N_noxref_15_1 0.00192258f
x_PM_AOI221xp5_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_AOI221xp5_ASAP7_75t_R%noxref_15
cc_66 N_noxref_15_1 N_MM0_g 0.00372181f
cc_67 N_noxref_15_1 N_NET012_8 0.000735421f
x_PM_AOI221xp5_ASAP7_75t_R%NET012 VSS N_MM1_d N_MM29_d N_MM31_d N_NET012_7
+ N_NET012_1 N_NET012_9 N_NET012_8 N_NET012_2 PM_AOI221xp5_ASAP7_75t_R%NET012
cc_68 N_NET012_7 N_C_1 0.000688371f
cc_69 N_NET012_1 N_C_4 0.000796799f
cc_70 N_NET012_1 N_MM28_g 0.000913798f
cc_71 N_NET012_7 N_MM28_g 0.0346771f
cc_72 N_NET012_7 N_A1_1 0.000780868f
cc_73 N_NET012_1 N_MM2_g 0.000896158f
cc_74 N_NET012_9 N_A1_4 0.0011027f
cc_75 N_NET012_1 N_A1_4 0.00132831f
cc_76 N_NET012_7 N_MM2_g 0.0342104f
cc_77 N_NET012_8 N_A2_1 0.000927448f
cc_78 N_NET012_2 N_MM0_g 0.00112538f
cc_79 N_NET012_9 N_A2_4 0.00134075f
cc_80 N_NET012_2 N_A2_4 0.00158618f
cc_81 N_NET012_8 N_MM0_g 0.0344957f
cc_82 N_NET012_7 N_NET16_8 0.000561226f
cc_83 N_NET012_9 N_NET16_9 0.00113994f
cc_84 N_NET012_1 N_NET16_2 0.00401665f
*END of AOI221xp5_ASAP7_75t_R.pxi
.ENDS
** Design:	AOI222xp33_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AOI222xp33_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AOI222xp33_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AOI222xp33_ASAP7_75t_R%NET49 VSS 2 3 1
c1 1 VSS 0.000851039f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0540 $X2=0.1080 $Y2=0.0540
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0540 $X2=0.1080 $Y2=0.0540
.ends

.subckt PM_AOI222xp33_ASAP7_75t_R%NET51 VSS 2 3 1
c1 1 VSS 0.000841852f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0540 $X2=0.2160 $Y2=0.0540
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0540 $X2=0.2160 $Y2=0.0540
.ends

.subckt PM_AOI222xp33_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.0425386f
.ends

.subckt PM_AOI222xp33_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.0328157f
.ends

.subckt PM_AOI222xp33_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.00640368f
.ends

.subckt PM_AOI222xp33_ASAP7_75t_R%NET50 VSS 2 3 1
c1 1 VSS 0.000857803f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0540 $X2=0.4320 $Y2=0.0540
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0540 $X2=0.4320 $Y2=0.0540
.ends

.subckt PM_AOI222xp33_ASAP7_75t_R%C2 VSS 8 3 1 4
c1 1 VSS 0.00359429f
c2 3 VSS 0.0717671f
c3 4 VSS 0.0173726f
r1 8 7 0.408082 $w=1.3e-08 $l=1.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1470 $X2=0.4590 $Y2=0.1452
r2 6 7 2.3902 $w=1.3e-08 $l=1.02e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1452
r3 4 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0980 $X2=0.4590 $Y2=0.1350
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r5 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1350
+ $X2=0.4590 $Y2=0.1350
.ends

.subckt PM_AOI222xp33_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.0417771f
.ends

.subckt PM_AOI222xp33_ASAP7_75t_R%NET27 VSS 16 17 31 32 7 1 9 8 11 2
c1 1 VSS 0.00328008f
c2 2 VSS 0.00976275f
c3 7 VSS 0.00239661f
c4 8 VSS 0.00481847f
c5 9 VSS 0.0030771f
c6 10 VSS 0.000826625f
c7 11 VSS 0.0113358f
c8 12 VSS 0.000914974f
c9 13 VSS 0.00297231f
r1 32 30 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r2 1 30 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r3 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r4 31 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r5 1 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.1980
r6 27 28 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1980 $X2=0.2295 $Y2=0.1980
r7 25 28 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1980 $X2=0.2295 $Y2=0.1980
r8 24 25 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2680
+ $Y=0.1980 $X2=0.2430 $Y2=0.1980
r9 9 12 7.11966 $w=1.35385e-08 $l=3.8396e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3130 $Y=0.1980 $X2=0.3510 $Y2=0.2035
r10 9 24 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3130
+ $Y=0.1980 $X2=0.2680 $Y2=0.1980
r11 10 13 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.2160 $X2=0.3510 $Y2=0.2340
r12 10 12 2.45586 $w=1.44e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.2160 $X2=0.3510 $Y2=0.2035
r13 13 21 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.2340 $X2=0.3780 $Y2=0.2340
r14 20 21 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r15 11 18 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4185
+ $Y=0.2340 $X2=0.4320 $Y2=0.2340
r16 11 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4185
+ $Y=0.2340 $X2=0.4050 $Y2=0.2340
r17 2 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.2340
r18 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r19 2 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r20 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r21 16 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
.ends

.subckt PM_AOI222xp33_ASAP7_75t_R%C1 VSS 6 3 1 4
c1 1 VSS 0.00657227f
c2 3 VSS 0.0461795f
c3 4 VSS 0.0055079f
r1 7 8 5.77145 $w=1.3e-08 $l=2.48e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1102 $X2=0.4050 $Y2=0.1350
r2 6 7 3.78933 $w=1.3e-08 $l=1.62e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0940 $X2=0.4050 $Y2=0.1102
r3 6 4 2.85657 $w=1.3e-08 $l=1.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0940 $X2=0.4050 $Y2=0.0817
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
.ends

.subckt PM_AOI222xp33_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00464992f
.ends

.subckt PM_AOI222xp33_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.0056075f
.ends

.subckt PM_AOI222xp33_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.00497817f
.ends

.subckt PM_AOI222xp33_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.00455485f
.ends

.subckt PM_AOI222xp33_ASAP7_75t_R%NET53 VSS 15 30 31 33 10 1 2 11 12 3 13
c1 1 VSS 0.00528824f
c2 2 VSS 0.00429579f
c3 3 VSS 0.00548053f
c4 10 VSS 0.00222182f
c5 11 VSS 0.00205431f
c6 12 VSS 0.00240171f
c7 13 VSS 0.0201801f
r1 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2680 $Y2=0.2025
r2 33 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r3 31 29 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r4 2 29 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r5 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r6 30 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r7 3 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.2340
r8 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r9 25 26 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2315
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r10 24 25 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2000
+ $Y=0.2340 $X2=0.2315 $Y2=0.2340
r11 23 24 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.2000 $Y2=0.2340
r12 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1755
+ $Y=0.2340 $X2=0.1890 $Y2=0.2340
r13 21 22 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r14 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r15 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1485 $Y2=0.2340
r16 18 19 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1240
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r17 17 18 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0925
+ $Y=0.2340 $X2=0.1240 $Y2=0.2340
r18 16 17 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2340 $X2=0.0925 $Y2=0.2340
r19 13 16 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r20 1 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r21 15 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r22 10 14 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r23 1 10 1e-05
.ends

.subckt PM_AOI222xp33_ASAP7_75t_R%A2 VSS 6 3 1 4
c1 1 VSS 0.00564293f
c2 3 VSS 0.0354533f
c3 4 VSS 0.00421698f
r1 7 8 4.37231 $w=1.3e-08 $l=1.88e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1162 $X2=0.1350 $Y2=0.1350
r2 6 7 2.39019 $w=1.3e-08 $l=1.02e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1060 $X2=0.1350 $Y2=0.1162
r3 6 4 4.25571 $w=1.3e-08 $l=1.83e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1060 $X2=0.1350 $Y2=0.0877
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AOI222xp33_ASAP7_75t_R%A1 VSS 8 3 1 4
c1 1 VSS 0.00649875f
c2 3 VSS 0.00843244f
c3 4 VSS 0.00414408f
r1 8 7 0.408082 $w=1.3e-08 $l=1.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1470 $X2=0.0810 $Y2=0.1452
r2 6 7 2.39019 $w=1.3e-08 $l=1.02e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1452
r3 4 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0980 $X2=0.0810 $Y2=0.1350
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r5 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AOI222xp33_ASAP7_75t_R%B2 VSS 8 3 1 4
c1 1 VSS 0.00601676f
c2 3 VSS 0.0355911f
c3 4 VSS 0.00423364f
r1 8 7 0.874462 $w=1.3e-08 $l=3.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1510 $X2=0.1890 $Y2=0.1472
r2 6 7 2.85657 $w=1.3e-08 $l=1.22e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1472
r3 4 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0980 $X2=0.1890 $Y2=0.1350
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r5 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AOI222xp33_ASAP7_75t_R%B1 VSS 6 3 1 4
c1 1 VSS 0.00700086f
c2 3 VSS 0.00905724f
c3 4 VSS 0.00493203f
r1 7 8 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1122 $X2=0.2430 $Y2=0.1350
r2 6 7 3.32295 $w=1.3e-08 $l=1.42e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0980 $X2=0.2430 $Y2=0.1122
r3 6 4 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0980 $X2=0.2430 $Y2=0.0837
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AOI222xp33_ASAP7_75t_R%Y VSS 43 23 47 49 57 58 2 1 19 18 16 13 17 14
+ 3 4 15 21
c1 1 VSS 0.00553515f
c2 2 VSS 0.00280447f
c3 3 VSS 0.00596647f
c4 4 VSS 0.00662396f
c5 13 VSS 0.0025881f
c6 14 VSS 0.00272797f
c7 15 VSS 0.00307487f
c8 16 VSS 0.00215547f
c9 17 VSS 0.00214274f
c10 18 VSS 0.0344046f
c11 19 VSS 0.000782942f
c12 20 VSS 0.00279706f
c13 21 VSS 0.000786815f
r1 58 56 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r2 2 56 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r3 16 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r4 57 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
r5 2 53 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.1980
r6 52 53 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.1980 $X2=0.1080 $Y2=0.1980
r7 51 52 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1980 $X2=0.0945 $Y2=0.1980
r8 50 51 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.0560
+ $Y=0.1980 $X2=0.0810 $Y2=0.1980
r9 19 21 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0380 $Y=0.1980 $X2=0.0270 $Y2=0.1980
r10 19 50 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0380
+ $Y=0.1980 $X2=0.0560 $Y2=0.1980
r11 21 45 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1980 $X2=0.0270 $Y2=0.1765
r12 49 48 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0540 $X2=0.3925 $Y2=0.0540
r13 15 48 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3800 $Y=0.0540 $X2=0.3925 $Y2=0.0540
r14 14 3 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0540 $X2=0.2680 $Y2=0.0540
r15 47 14 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0540 $X2=0.2555 $Y2=0.0540
r16 44 45 4.83869 $w=1.3e-08 $l=2.08e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1557 $X2=0.0270 $Y2=0.1765
r17 43 44 2.04041 $w=1.3e-08 $l=8.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1470 $X2=0.0270 $Y2=0.1557
r18 43 42 9.0361 $w=1.3e-08 $l=3.88e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1470 $X2=0.0270 $Y2=0.1082
r19 17 20 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0575 $X2=0.0270 $Y2=0.0360
r20 17 42 11.8344 $w=1.3e-08 $l=5.07e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0575 $X2=0.0270 $Y2=0.1082
r21 4 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.0540
+ $X2=0.3780 $Y2=0.0360
r22 3 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0540
+ $X2=0.2700 $Y2=0.0360
r23 38 39 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3645
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r24 37 38 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3195
+ $Y=0.0360 $X2=0.3645 $Y2=0.0360
r25 36 37 11.5429 $w=1.3e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.3195 $Y2=0.0360
r26 35 36 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r27 34 35 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2565 $Y2=0.0360
r28 33 34 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2180
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r29 32 33 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2000
+ $Y=0.0360 $X2=0.2180 $Y2=0.0360
r30 31 32 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.2000 $Y2=0.0360
r31 30 31 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r32 29 30 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r33 28 29 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1240
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r34 27 28 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1060
+ $Y=0.0360 $X2=0.1240 $Y2=0.0360
r35 26 27 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0360 $X2=0.1060 $Y2=0.0360
r36 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0675
+ $Y=0.0360 $X2=0.0810 $Y2=0.0360
r37 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.0360 $X2=0.0675 $Y2=0.0360
r38 18 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r39 18 20 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0405 $Y=0.0360 $X2=0.0270 $Y2=0.0360
r40 1 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0540 $Y2=0.0360
r41 23 22 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r42 13 22 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r43 4 15 1e-05
r44 1 13 1e-05
.ends


*
.SUBCKT AOI222xp33_ASAP7_75t_R VSS VDD A1 A2 B2 B1 C1 C2 Y
*
* VSS VSS
* VDD VDD
* A1 A1
* A2 A2
* B2 B2
* B1 B1
* C1 C1
* C2 C2
* Y Y
*
*

MM0 N_MM0_d N_MM0_g N_MM0_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1 N_MM1_d N_MM1_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM4 N_MM4_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g N_MM3_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM7_g N_MM5_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM6 N_MM6_d N_MM10_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM9 N_MM9_d N_MM0_g N_MM9_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM12 N_MM12_d N_MM1_g N_MM12_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 N_MM11_d N_MM4_g N_MM11_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM3_g N_MM8_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AOI222xp33_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AOI222xp33_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AOI222xp33_ASAP7_75t_R%NET49 VSS N_MM0_s N_MM1_d N_NET49_1
+ PM_AOI222xp33_ASAP7_75t_R%NET49
cc_1 N_NET49_1 N_MM0_g 0.012498f
cc_2 N_NET49_1 N_MM1_g 0.0125363f
x_PM_AOI222xp33_ASAP7_75t_R%NET51 VSS N_MM4_d N_MM3_s N_NET51_1
+ PM_AOI222xp33_ASAP7_75t_R%NET51
cc_3 N_NET51_1 N_MM4_g 0.0126497f
cc_4 N_NET51_1 N_MM3_g 0.0127291f
x_PM_AOI222xp33_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_AOI222xp33_ASAP7_75t_R%noxref_22
cc_5 N_noxref_22_1 N_MM10_g 0.00182863f
cc_6 N_noxref_22_1 N_noxref_21_1 0.00192757f
x_PM_AOI222xp33_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_AOI222xp33_ASAP7_75t_R%noxref_21
cc_7 N_noxref_21_1 N_MM10_g 0.00378185f
x_PM_AOI222xp33_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_AOI222xp33_ASAP7_75t_R%noxref_18
cc_8 N_noxref_18_1 N_MM3_g 0.00151756f
cc_9 N_noxref_18_1 N_NET53_12 0.0360402f
cc_10 N_noxref_18_1 N_noxref_17_1 0.00133951f
x_PM_AOI222xp33_ASAP7_75t_R%NET50 VSS N_MM5_s N_MM6_d N_NET50_1
+ PM_AOI222xp33_ASAP7_75t_R%NET50
cc_11 N_NET50_1 N_MM7_g 0.012587f
cc_12 N_NET50_1 N_MM10_g 0.0126504f
x_PM_AOI222xp33_ASAP7_75t_R%C2 VSS C2 N_MM10_g N_C2_1 N_C2_4
+ PM_AOI222xp33_ASAP7_75t_R%C2
cc_13 N_C2_1 N_C1_1 0.00137255f
cc_14 N_C2_4 N_C1_4 0.0055703f
cc_15 N_MM10_g N_MM7_g 0.00773099f
x_PM_AOI222xp33_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_AOI222xp33_ASAP7_75t_R%noxref_20
cc_16 N_noxref_20_1 N_MM7_g 0.00154311f
cc_17 N_noxref_20_1 N_NET53_12 0.000541884f
cc_18 N_noxref_20_1 N_noxref_17_1 0.000475614f
cc_19 N_noxref_20_1 N_noxref_18_1 0.00764323f
cc_20 N_noxref_20_1 N_noxref_19_1 0.00135354f
x_PM_AOI222xp33_ASAP7_75t_R%NET27 VSS N_MM7_d N_MM10_d N_MM11_s N_MM8_s
+ N_NET27_7 N_NET27_1 N_NET27_9 N_NET27_8 N_NET27_11 N_NET27_2
+ PM_AOI222xp33_ASAP7_75t_R%NET27
cc_21 N_NET27_7 N_B2_4 0.000575605f
cc_22 N_NET27_1 N_B2_4 0.000771546f
cc_23 N_NET27_7 N_B2_1 0.000780398f
cc_24 N_NET27_1 N_MM4_g 0.000891671f
cc_25 N_NET27_7 N_MM4_g 0.0339735f
cc_26 N_NET27_7 N_B1_1 0.000826548f
cc_27 N_NET27_1 N_MM3_g 0.000896182f
cc_28 N_NET27_9 N_B1_4 0.00140103f
cc_29 N_NET27_1 N_B1_4 0.00152652f
cc_30 N_NET27_7 N_MM3_g 0.0341573f
cc_31 N_NET27_8 N_C1_4 0.000538813f
cc_32 N_NET27_8 N_C1_1 0.000608449f
cc_33 N_NET27_11 N_C1_4 0.00108431f
cc_34 N_NET27_2 N_MM7_g 0.00117987f
cc_35 N_NET27_2 N_C1_4 0.00226075f
cc_36 N_NET27_8 N_MM7_g 0.0345444f
cc_37 N_NET27_11 N_C2_4 0.000960587f
cc_38 N_NET27_2 N_MM10_g 0.00120663f
cc_39 N_NET27_2 N_C2_4 0.00156893f
cc_40 N_NET27_8 N_MM10_g 0.0346646f
cc_41 N_NET27_9 N_NET53_11 0.000561689f
cc_42 N_NET27_7 N_NET53_12 0.00175569f
cc_43 N_NET27_1 N_NET53_13 0.000777485f
cc_44 N_NET27_1 N_NET53_2 0.0013397f
cc_45 N_NET27_1 N_NET53_3 0.00498503f
cc_46 N_NET27_9 N_NET53_13 0.0100124f
x_PM_AOI222xp33_ASAP7_75t_R%C1 VSS C1 N_MM7_g N_C1_1 N_C1_4
+ PM_AOI222xp33_ASAP7_75t_R%C1
x_PM_AOI222xp33_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_AOI222xp33_ASAP7_75t_R%noxref_15
cc_47 N_noxref_15_1 N_MM0_g 0.00350361f
cc_48 N_noxref_15_1 N_Y_1 0.000430399f
cc_49 N_noxref_15_1 N_Y_13 0.027578f
cc_50 N_noxref_15_1 N_NET53_10 0.000580839f
x_PM_AOI222xp33_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_AOI222xp33_ASAP7_75t_R%noxref_16
cc_51 N_noxref_16_1 N_MM0_g 0.00159707f
cc_52 N_noxref_16_1 N_Y_16 0.000872388f
cc_53 N_noxref_16_1 N_NET53_10 0.0363942f
cc_54 N_noxref_16_1 N_noxref_15_1 0.0019015f
x_PM_AOI222xp33_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_AOI222xp33_ASAP7_75t_R%noxref_19
cc_55 N_noxref_19_1 N_MM7_g 0.00345578f
cc_56 N_noxref_19_1 N_Y_15 0.0276018f
cc_57 N_noxref_19_1 N_noxref_17_1 0.00777986f
cc_58 N_noxref_19_1 N_noxref_18_1 0.00046902f
x_PM_AOI222xp33_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_AOI222xp33_ASAP7_75t_R%noxref_17
cc_59 N_noxref_17_1 N_MM3_g 0.00344651f
cc_60 N_noxref_17_1 N_Y_14 0.0276002f
cc_61 N_noxref_17_1 N_NET53_12 0.000479905f
x_PM_AOI222xp33_ASAP7_75t_R%NET53 VSS N_MM9_s N_MM12_s N_MM11_d N_MM8_d
+ N_NET53_10 N_NET53_1 N_NET53_2 N_NET53_11 N_NET53_12 N_NET53_3 N_NET53_13
+ PM_AOI222xp33_ASAP7_75t_R%NET53
cc_62 N_NET53_10 N_A1_1 0.000855343f
cc_63 N_NET53_1 N_MM0_g 0.00103719f
cc_64 N_NET53_10 N_MM0_g 0.0345609f
cc_65 N_NET53_2 N_MM1_g 0.00142938f
cc_66 N_NET53_11 N_A2_1 0.000779372f
cc_67 N_NET53_11 N_MM1_g 0.0342612f
cc_68 N_NET53_11 N_B2_1 0.000775665f
cc_69 N_NET53_2 N_MM4_g 0.000982368f
cc_70 N_NET53_11 N_MM4_g 0.0347075f
cc_71 N_NET53_12 N_B1_1 0.000870848f
cc_72 N_NET53_3 N_MM3_g 0.00112691f
cc_73 N_NET53_12 N_MM3_g 0.0348528f
cc_74 N_NET53_13 N_Y_16 0.000564156f
cc_75 N_NET53_13 N_Y_21 0.000632052f
cc_76 N_NET53_10 N_Y_16 0.000712084f
cc_77 N_NET53_1 N_Y_17 0.000726767f
cc_78 N_NET53_1 N_Y_19 0.000775922f
cc_79 N_NET53_13 N_Y_2 0.000792769f
cc_80 N_NET53_11 N_Y_16 0.0011243f
cc_81 N_NET53_1 N_Y_2 0.00240982f
cc_82 N_NET53_2 N_Y_2 0.00417564f
cc_83 N_NET53_13 N_Y_19 0.00866358f
x_PM_AOI222xp33_ASAP7_75t_R%A2 VSS A2 N_MM1_g N_A2_1 N_A2_4
+ PM_AOI222xp33_ASAP7_75t_R%A2
cc_84 N_A2_1 N_A1_1 0.00131028f
cc_85 N_A2_4 N_A1_4 0.00339487f
cc_86 N_MM1_g N_MM0_g 0.00756334f
x_PM_AOI222xp33_ASAP7_75t_R%A1 VSS A1 N_MM0_g N_A1_1 N_A1_4
+ PM_AOI222xp33_ASAP7_75t_R%A1
x_PM_AOI222xp33_ASAP7_75t_R%B2 VSS B2 N_MM4_g N_B2_1 N_B2_4
+ PM_AOI222xp33_ASAP7_75t_R%B2
cc_87 N_B2_1 N_A2_1 0.00129724f
cc_88 N_B2_4 N_A2_4 0.00338386f
cc_89 N_MM4_g N_MM1_g 0.00635668f
x_PM_AOI222xp33_ASAP7_75t_R%B1 VSS B1 N_MM3_g N_B1_1 N_B1_4
+ PM_AOI222xp33_ASAP7_75t_R%B1
cc_90 N_B1_1 N_B2_1 0.00138836f
cc_91 N_B1_4 N_B2_4 0.00365367f
cc_92 N_MM3_g N_MM4_g 0.00757174f
x_PM_AOI222xp33_ASAP7_75t_R%Y VSS Y N_MM0_d N_MM3_d N_MM5_d N_MM9_d N_MM12_d
+ N_Y_2 N_Y_1 N_Y_19 N_Y_18 N_Y_16 N_Y_13 N_Y_17 N_Y_14 N_Y_3 N_Y_4 N_Y_15
+ N_Y_21 PM_AOI222xp33_ASAP7_75t_R%Y
cc_93 N_Y_2 N_A1_1 0.000766015f
cc_94 N_Y_2 N_MM0_g 0.000919422f
cc_95 N_Y_1 N_MM0_g 0.000938199f
cc_96 N_Y_19 N_A1_4 0.00111274f
cc_97 N_Y_18 N_A1_4 0.00122712f
cc_98 N_Y_16 N_A1_1 0.00132923f
cc_99 N_Y_13 N_MM0_g 0.0108411f
cc_100 N_Y_17 N_A1_4 0.00661683f
cc_101 N_Y_16 N_MM0_g 0.0492846f
cc_102 N_Y_2 N_MM1_g 0.00127011f
cc_103 N_Y_19 N_A2_4 0.000552156f
cc_104 N_Y_16 N_A2_1 0.000881115f
cc_105 N_Y_18 N_A2_4 0.001376f
cc_106 N_Y_2 N_A2_4 0.00219552f
cc_107 N_Y_16 N_MM1_g 0.03537f
cc_108 N_Y_16 N_B2_4 0.000270598f
cc_109 N_Y_18 N_B2_4 0.00353933f
cc_110 N_Y_14 N_B1_1 0.000397068f
cc_111 N_Y_3 N_MM3_g 0.00105247f
cc_112 N_Y_18 N_B1_4 0.00165515f
cc_113 N_Y_3 N_B1_4 0.00212848f
cc_114 N_Y_14 N_MM3_g 0.0258012f
cc_115 N_Y_18 N_C1_4 0.0010492f
cc_116 N_Y_4 N_MM7_g 0.00107847f
cc_117 N_Y_4 N_C1_4 0.00158291f
cc_118 N_Y_15 N_MM7_g 0.0259866f
*END of AOI222xp33_ASAP7_75t_R.pxi
.ENDS
** Design:	AOI22x1_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AOI22x1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AOI22x1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AOI22x1_ASAP7_75t_R%NET30__2 VSS 2 3 1
c1 1 VSS 0.0009531f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3240 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3240 $Y2=0.0675
.ends

.subckt PM_AOI22x1_ASAP7_75t_R%NET30 VSS 2 3 1
c1 1 VSS 0.000970173f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4320 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4320 $Y2=0.0675
.ends

.subckt PM_AOI22x1_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.011557f
.ends

.subckt PM_AOI22x1_ASAP7_75t_R%A1 VSS 21 3 4 6 1 7
c1 1 VSS 0.0116502f
c2 3 VSS 0.0468451f
c3 4 VSS 0.0469385f
c4 5 VSS 0.00355196f
c5 6 VSS 0.00420478f
c6 7 VSS 0.00349407f
r1 21 22 0.0765333 $w=1.8e-08 $l=7e-10 $layer=M1 $thickness=3.6e-08 $X=0.3590
+ $Y=0.1620 $X2=0.3597 $Y2=0.1620
r2 21 7 0.892889 $w=1.8e-08 $l=8.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.3590
+ $Y=0.1620 $X2=0.3502 $Y2=0.1620
r3 7 18 0.958461 $w=1.77143e-08 $l=9.53362e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.3502 $Y=0.1620 $X2=0.3510 $Y2=0.1525
r4 4 16 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r5 18 22 0.142106 $w=1.46667e-08 $l=1.28818e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.1525 $X2=0.3597 $Y2=0.1620
r6 5 9 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1345
+ $X2=0.3510 $Y2=0.1350
r7 5 18 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1345 $X2=0.3510 $Y2=0.1525
r8 5 6 4.99922 $w=1.46981e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.1345 $X2=0.3510 $Y2=0.1080
r9 14 16 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3925 $Y=0.1350 $X2=0.4050 $Y2=0.1350
r10 13 14 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3780 $Y=0.1350 $X2=0.3925 $Y2=0.1350
r11 12 13 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3635 $Y=0.1350 $X2=0.3780 $Y2=0.1350
r12 10 12 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.3605 $Y=0.1350 $X2=0.3635 $Y2=0.1350
r13 9 10 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3605 $Y2=0.1350
r14 1 9 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.3415
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r15 1 11 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.3415
+ $Y=0.1350 $X2=0.3405 $Y2=0.1350
r16 3 9 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r17 3 11 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.3510 $Y=0.1350 $X2=0.3405 $Y2=0.1350
r18 3 12 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.3510 $Y=0.1350 $X2=0.3635 $Y2=0.1350
.ends

.subckt PM_AOI22x1_ASAP7_75t_R%NET29__2 VSS 2 3 1
c1 1 VSS 0.000961773f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_AOI22x1_ASAP7_75t_R%NET29 VSS 2 3 1
c1 1 VSS 0.000954862f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2160 $Y2=0.0675
.ends

.subckt PM_AOI22x1_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00577845f
.ends

.subckt PM_AOI22x1_ASAP7_75t_R%B1 VSS 23 3 4 6 5 1 7
c1 1 VSS 0.0136717f
c2 3 VSS 0.0843442f
c3 4 VSS 0.0844316f
c4 5 VSS 0.00340528f
c5 6 VSS 0.00359845f
c6 7 VSS 0.00313732f
r1 7 21 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1980 $X2=0.1890 $Y2=0.1800
r2 23 24 0.790844 $w=1.8e-08 $l=7.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1830
+ $Y=0.1080 $X2=0.1907 $Y2=0.1080
r3 23 6 0.178578 $w=1.8e-08 $l=1.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.1830
+ $Y=0.1080 $X2=0.1812 $Y2=0.1080
r4 3 15 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r5 20 21 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1625 $X2=0.1890 $Y2=0.1800
r6 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1490 $X2=0.1890 $Y2=0.1625
r7 18 19 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1490
r8 5 18 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1215 $X2=0.1890 $Y2=0.1350
r9 5 24 1.78918 $w=1.60851e-08 $l=1.36066e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1215 $X2=0.1907 $Y2=0.1080
r10 13 15 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1475 $Y=0.1350 $X2=0.1350 $Y2=0.1350
r11 12 13 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1620 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r12 11 12 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1765 $Y=0.1350 $X2=0.1620 $Y2=0.1350
r13 10 17 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1985 $Y=0.1350 $X2=0.1995 $Y2=0.1350
r14 9 10 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1985 $Y2=0.1350
r15 9 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
r16 1 9 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1795
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r17 1 11 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1795 $Y=0.1350 $X2=0.1765 $Y2=0.1350
r18 4 9 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r19 4 11 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1765 $Y2=0.1350
r20 4 17 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.1890 $Y=0.1350 $X2=0.1995 $Y2=0.1350
.ends

.subckt PM_AOI22x1_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00626074f
.ends

.subckt PM_AOI22x1_ASAP7_75t_R%A2 VSS 20 5 6 10 7 1 8 2 12 9 11
c1 1 VSS 0.00556892f
c2 2 VSS 0.00549685f
c3 5 VSS 0.00811502f
c4 6 VSS 0.00779892f
c5 7 VSS 0.00339354f
c6 8 VSS 0.00585128f
c7 9 VSS 0.00310501f
c8 10 VSS 0.00291221f
c9 11 VSS 0.00285482f
c10 12 VSS 0.00290142f
r1 2 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1350
+ $X2=0.4590 $Y2=0.1350
r2 6 2 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r3 11 29 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1620 $X2=0.4590 $Y2=0.1485
r4 28 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1485
r5 27 28 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1215 $X2=0.4590 $Y2=0.1350
r6 26 27 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1080 $X2=0.4590 $Y2=0.1215
r7 9 12 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0900 $X2=0.4590 $Y2=0.0720
r8 9 26 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0900 $X2=0.4590 $Y2=0.1080
r9 12 25 2.6649 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0720 $X2=0.4405 $Y2=0.0720
r10 24 25 8.27824 $w=1.3e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0720 $X2=0.4405 $Y2=0.0720
r11 23 24 10.3769 $w=1.3e-08 $l=4.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3605
+ $Y=0.0720 $X2=0.4050 $Y2=0.0720
r12 22 23 8.16164 $w=1.3e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3255
+ $Y=0.0720 $X2=0.3605 $Y2=0.0720
r13 8 10 0.79938 $w=1.72857e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3075 $Y=0.0720 $X2=0.2970 $Y2=0.0720
r14 8 22 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3075
+ $Y=0.0720 $X2=0.3255 $Y2=0.0720
r15 10 19 1.09087 $w=2.05064e-08 $l=1.17e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0720 $X2=0.2970 $Y2=0.0837
r16 20 21 1.45744 $w=1.3e-08 $l=6.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0870 $X2=0.2970 $Y2=0.0932
r17 20 19 0.757867 $w=1.3e-08 $l=3.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0870 $X2=0.2970 $Y2=0.0837
r18 18 21 3.43955 $w=1.3e-08 $l=1.48e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1080 $X2=0.2970 $Y2=0.0932
r19 7 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1215 $X2=0.2970 $Y2=0.1350
r20 7 18 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1215 $X2=0.2970 $Y2=0.1080
r21 5 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r22 1 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_AOI22x1_ASAP7_75t_R%B2 VSS 18 5 6 7 2 9 1 8 12 11 10
c1 1 VSS 0.00617676f
c2 2 VSS 0.00625371f
c3 5 VSS 0.0451832f
c4 6 VSS 0.0453254f
c5 7 VSS 0.00382326f
c6 8 VSS 0.00531878f
c7 9 VSS 0.00301784f
c8 10 VSS 0.00241633f
c9 11 VSS 0.0035509f
c10 12 VSS 0.00231447f
r1 2 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
r2 6 2 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r3 27 28 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1215 $X2=0.2430 $Y2=0.1350
r4 26 27 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1080 $X2=0.2430 $Y2=0.1215
r5 9 12 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0900 $X2=0.2430 $Y2=0.0720
r6 9 26 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0900 $X2=0.2430 $Y2=0.1080
r7 12 25 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0720 $X2=0.2160 $Y2=0.0720
r8 24 25 8.51143 $w=1.3e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.1795
+ $Y=0.0720 $X2=0.2160 $Y2=0.0720
r9 23 24 10.3769 $w=1.3e-08 $l=4.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0720 $X2=0.1795 $Y2=0.0720
r10 8 10 2.6649 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0995 $Y=0.0720 $X2=0.0810 $Y2=0.0720
r11 8 23 8.27824 $w=1.3e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.0995
+ $Y=0.0720 $X2=0.1350 $Y2=0.0720
r12 11 21 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1980 $X2=0.0810 $Y2=0.1665
r13 10 16 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0720 $X2=0.0810 $Y2=0.0900
r14 20 21 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1665
r15 19 20 2.97317 $w=1.3e-08 $l=1.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1222 $X2=0.0810 $Y2=0.1350
r16 18 19 0.991057 $w=1.3e-08 $l=4.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1180 $X2=0.0810 $Y2=0.1222
r17 18 17 0.174892 $w=1.3e-08 $l=8e-10 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1180 $X2=0.0810 $Y2=0.1172
r18 7 16 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1080 $X2=0.0810 $Y2=0.0900
r19 7 17 2.15701 $w=1.3e-08 $l=9.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1080 $X2=0.0810 $Y2=0.1172
r20 5 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r21 1 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AOI22x1_ASAP7_75t_R%NET13 VSS 24 25 46 49 50 53 54 56 18 3 16 1 21 2
+ 17 20 5 4 19
c1 1 VSS 0.00802004f
c2 2 VSS 0.00972443f
c3 3 VSS 0.007137f
c4 4 VSS 0.00417834f
c5 5 VSS 0.00521762f
c6 16 VSS 0.00343005f
c7 17 VSS 0.00446098f
c8 18 VSS 0.00321387f
c9 19 VSS 0.00206973f
c10 20 VSS 0.00220256f
c11 21 VSS 0.0383791f
r1 20 5 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4840 $Y2=0.2025
r2 56 20 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r3 54 52 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r4 4 52 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r5 19 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3780 $Y2=0.2025
r6 53 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r7 50 48 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r8 3 48 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r9 18 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r10 49 18 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r11 46 45 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r12 16 45 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r13 5 43 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2025
+ $X2=0.4860 $Y2=0.2340
r14 4 41 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.2340
r15 3 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.2340
r16 1 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r17 42 43 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4860 $Y2=0.2340
r18 41 42 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.4320 $Y2=0.2340
r19 40 41 9.0944 $w=1.3e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.3390
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r20 39 40 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3075
+ $Y=0.2340 $X2=0.3390 $Y2=0.2340
r21 38 39 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.2340 $X2=0.3075 $Y2=0.2340
r22 37 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2835
+ $Y=0.2340 $X2=0.2970 $Y2=0.2340
r23 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.2835 $Y2=0.2340
r24 35 36 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r25 34 35 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2565 $Y2=0.2340
r26 33 34 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2430 $Y2=0.2340
r27 32 33 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1845
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r28 31 32 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1660
+ $Y=0.2340 $X2=0.1845 $Y2=0.2340
r29 29 30 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2340 $X2=0.0675 $Y2=0.2340
r30 27 30 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.0905
+ $Y=0.2340 $X2=0.0675 $Y2=0.2340
r31 26 31 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1570
+ $Y=0.2340 $X2=0.1660 $Y2=0.2340
r32 21 26 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.1310
+ $Y=0.2340 $X2=0.1570 $Y2=0.2340
r33 21 27 9.44418 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1310
+ $Y=0.2340 $X2=0.0905 $Y2=0.2340
r34 2 31 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1660 $Y2=0.2340
r35 24 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r36 2 23 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r37 17 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r38 25 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r39 1 16 1e-05
.ends

.subckt PM_AOI22x1_ASAP7_75t_R%Y VSS 44 27 41 42 49 61 62 65 66 1 17 2 16 21 20
+ 19 3 4 5 23 22 18 25
c1 1 VSS 0.00621494f
c2 2 VSS 0.00556792f
c3 3 VSS 0.00290372f
c4 4 VSS 0.00282979f
c5 5 VSS 0.00573507f
c6 16 VSS 0.0032369f
c7 17 VSS 0.00320621f
c8 18 VSS 0.00266664f
c9 19 VSS 0.0021207f
c10 20 VSS 0.00210863f
c11 21 VSS 0.0428987f
c12 22 VSS 0.00143258f
c13 23 VSS 0.00205739f
c14 24 VSS 0.00273476f
c15 25 VSS 0.000747503f
r1 66 64 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r2 3 64 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r3 19 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r4 65 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r5 62 60 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r6 4 60 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r7 20 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r8 61 20 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r9 3 57 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.1980
r10 4 51 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4360 $Y2=0.1980
r11 57 58 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1980 $X2=0.3375 $Y2=0.1980
r12 55 58 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.3605
+ $Y=0.1980 $X2=0.3375 $Y2=0.1980
r13 53 54 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.4010
+ $Y=0.1980 $X2=0.4270 $Y2=0.1980
r14 53 55 9.44418 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4010
+ $Y=0.1980 $X2=0.3605 $Y2=0.1980
r15 51 52 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4360
+ $Y=0.1980 $X2=0.4545 $Y2=0.1980
r16 51 54 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4360
+ $Y=0.1980 $X2=0.4270 $Y2=0.1980
r17 50 52 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4840
+ $Y=0.1980 $X2=0.4545 $Y2=0.1980
r18 22 25 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5020 $Y=0.1980 $X2=0.5130 $Y2=0.1980
r19 22 50 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5020
+ $Y=0.1980 $X2=0.4840 $Y2=0.1980
r20 25 47 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1980 $X2=0.5130 $Y2=0.1800
r21 18 5 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0675 $X2=0.4840 $Y2=0.0675
r22 49 18 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4715 $Y2=0.0675
r23 46 47 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1620 $X2=0.5130 $Y2=0.1800
r24 45 46 6.58761 $w=1.3e-08 $l=2.83e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1337 $X2=0.5130 $Y2=0.1620
r25 44 45 4.6055 $w=1.3e-08 $l=1.97e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1140 $X2=0.5130 $Y2=0.1337
r26 44 43 6.00464 $w=1.3e-08 $l=2.58e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1140 $X2=0.5130 $Y2=0.0882
r27 23 24 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0540 $X2=0.5130 $Y2=0.0360
r28 23 43 7.98675 $w=1.3e-08 $l=3.42e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0540 $X2=0.5130 $Y2=0.0882
r29 42 40 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r30 2 40 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r31 17 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r32 41 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
r33 5 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0675
+ $X2=0.4860 $Y2=0.0360
r34 24 38 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.0360 $X2=0.4995 $Y2=0.0360
r35 2 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2700 $Y2=0.0360
r36 37 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.0360 $X2=0.4995 $Y2=0.0360
r37 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4725
+ $Y=0.0360 $X2=0.4860 $Y2=0.0360
r38 35 36 22.0364 $w=1.3e-08 $l=9.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0360 $X2=0.4725 $Y2=0.0360
r39 34 35 22.0364 $w=1.3e-08 $l=9.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.2835
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r40 33 34 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.2835 $Y2=0.0360
r41 32 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r42 31 32 22.0364 $w=1.3e-08 $l=9.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.2565 $Y2=0.0360
r43 30 31 22.0364 $w=1.3e-08 $l=9.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.0675
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r44 29 30 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.0360 $X2=0.0675 $Y2=0.0360
r45 28 29 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r46 21 28 0.816164 $w=1.3e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0390
+ $Y=0.0360 $X2=0.0425 $Y2=0.0360
r47 1 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0540 $Y2=0.0360
r48 27 26 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r49 16 26 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r50 1 16 1e-05
.ends


*
.SUBCKT AOI22x1_ASAP7_75t_R VSS VDD B2 B1 A2 A1 Y
*
* VSS VSS
* VDD VDD
* B2 B2
* B1 B1
* A2 A2
* A1 A1
* Y Y
*
*

MM7@2 N_MM7@2_d N_MM7@2_g N_MM7@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9@2 N_MM9@2_d N_MM9@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM2@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM3@2_g N_MM7_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6@2 N_MM6@2_d N_MM5_g N_MM6@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8@2 N_MM8@2_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM4@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM5@2_g N_MM6_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM7@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM9@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2@2 N_MM2@2_d N_MM2@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3@2 N_MM3@2_d N_MM3@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g N_MM4_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@2 N_MM4@2_d N_MM4@2_g N_MM4@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@2 N_MM5@2_d N_MM5@2_g N_MM5@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AOI22x1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AOI22x1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AOI22x1_ASAP7_75t_R%NET30__2 VSS N_MM6@2_s N_MM8@2_d N_NET30__2_1
+ PM_AOI22x1_ASAP7_75t_R%NET30__2
cc_1 N_NET30__2_1 N_MM5_g 0.017464f
cc_2 N_NET30__2_1 N_MM4_g 0.0174435f
x_PM_AOI22x1_ASAP7_75t_R%NET30 VSS N_MM8_d N_MM6_s N_NET30_1
+ PM_AOI22x1_ASAP7_75t_R%NET30
cc_3 N_NET30_1 N_MM5@2_g 0.0172989f
cc_4 N_NET30_1 N_MM4@2_g 0.0174847f
x_PM_AOI22x1_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_AOI22x1_ASAP7_75t_R%noxref_15
cc_5 N_noxref_15_1 N_MM5@2_g 0.00375941f
cc_6 N_noxref_15_1 N_NET13_20 0.0369825f
cc_7 N_noxref_15_1 N_Y_5 0.000616808f
cc_8 N_noxref_15_1 N_Y_18 0.0386863f
x_PM_AOI22x1_ASAP7_75t_R%A1 VSS A1 N_MM4_g N_MM4@2_g N_A1_6 N_A1_1 N_A1_7
+ PM_AOI22x1_ASAP7_75t_R%A1
cc_9 N_A1_6 N_A2_7 0.00197189f
cc_10 N_A1_1 N_A2_1 0.00341139f
cc_11 N_MM4@2_g N_MM5@2_g 0.00506948f
cc_12 N_MM4_g N_MM5_g 0.00507602f
cc_13 N_A1_6 N_A2_8 0.007793f
x_PM_AOI22x1_ASAP7_75t_R%NET29__2 VSS N_MM7@2_s N_MM9@2_d N_NET29__2_1
+ PM_AOI22x1_ASAP7_75t_R%NET29__2
cc_14 N_NET29__2_1 N_MM7@2_g 0.017261f
cc_15 N_NET29__2_1 N_MM9@2_g 0.0172581f
x_PM_AOI22x1_ASAP7_75t_R%NET29 VSS N_MM9_d N_MM7_s N_NET29_1
+ PM_AOI22x1_ASAP7_75t_R%NET29
cc_16 N_NET29_1 N_MM3@2_g 0.0173847f
cc_17 N_NET29_1 N_MM2@2_g 0.0175219f
x_PM_AOI22x1_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_AOI22x1_ASAP7_75t_R%noxref_13
cc_18 N_noxref_13_1 N_MM7@2_g 0.00165813f
cc_19 N_noxref_13_1 N_NET13_16 0.000555954f
cc_20 N_noxref_13_1 N_Y_16 0.0365586f
x_PM_AOI22x1_ASAP7_75t_R%B1 VSS B1 N_MM9@2_g N_MM2@2_g N_B1_6 N_B1_5 N_B1_1
+ N_B1_7 PM_AOI22x1_ASAP7_75t_R%B1
cc_21 N_B1_6 N_B2_7 0.00062908f
cc_22 N_B1_6 N_B2_2 0.00106522f
cc_23 N_B1_6 N_B2_9 0.00129672f
cc_24 N_B1_5 N_B2_9 0.00133753f
cc_25 N_B1_1 N_B2_1 0.00240154f
cc_26 N_MM9@2_g N_MM7@2_g 0.00507265f
cc_27 N_MM2@2_g N_MM3@2_g 0.00508937f
cc_28 N_B1_6 N_B2_8 0.00738468f
x_PM_AOI22x1_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_AOI22x1_ASAP7_75t_R%noxref_14
cc_29 N_noxref_14_1 N_MM7@2_g 0.00164466f
cc_30 N_noxref_14_1 N_NET13_16 0.0360749f
cc_31 N_noxref_14_1 N_Y_16 0.000566325f
cc_32 N_noxref_14_1 N_noxref_13_1 0.00179741f
x_PM_AOI22x1_ASAP7_75t_R%A2 VSS A2 N_MM5_g N_MM5@2_g N_A2_10 N_A2_7 N_A2_1
+ N_A2_8 N_A2_2 N_A2_12 N_A2_9 N_A2_11 PM_AOI22x1_ASAP7_75t_R%A2
cc_33 N_A2_10 N_B2_12 0.000845128f
cc_34 N_A2_7 N_B2_9 0.00283436f
cc_35 N_MM5_g N_MM3@2_g 0.00504601f
x_PM_AOI22x1_ASAP7_75t_R%B2 VSS B2 N_MM7@2_g N_MM3@2_g N_B2_7 N_B2_2 N_B2_9
+ N_B2_1 N_B2_8 N_B2_12 N_B2_11 N_B2_10 PM_AOI22x1_ASAP7_75t_R%B2
x_PM_AOI22x1_ASAP7_75t_R%NET13 VSS N_MM2@2_d N_MM2_d N_MM3_d N_MM3@2_d N_MM5_s
+ N_MM4_s N_MM4@2_s N_MM5@2_s N_NET13_18 N_NET13_3 N_NET13_16 N_NET13_1
+ N_NET13_21 N_NET13_2 N_NET13_17 N_NET13_20 N_NET13_5 N_NET13_4 N_NET13_19
+ PM_AOI22x1_ASAP7_75t_R%NET13
cc_36 N_NET13_18 N_MM3@2_g 0.0334448f
cc_37 N_NET13_3 N_B2_9 0.000429491f
cc_38 N_NET13_18 N_B2_2 0.000705419f
cc_39 N_NET13_16 N_B2_1 0.000755844f
cc_40 N_NET13_1 N_B2_7 0.000889737f
cc_41 N_NET13_3 N_MM3@2_g 0.00094434f
cc_42 N_NET13_1 N_MM7@2_g 0.00158106f
cc_43 N_NET13_21 N_B2_11 0.0023995f
cc_44 N_NET13_21 N_B2_9 0.00268879f
cc_45 N_NET13_16 N_MM7@2_g 0.0347908f
cc_46 N_NET13_2 N_MM9@2_g 0.00310134f
cc_47 N_NET13_17 N_B1_1 0.00243302f
cc_48 N_NET13_21 N_B1_7 0.0050239f
cc_49 N_NET13_17 N_MM2@2_g 0.018363f
cc_50 N_NET13_17 N_MM9@2_g 0.0497145f
cc_51 N_NET13_3 N_MM5_g 0.00122926f
cc_52 N_NET13_21 N_MM5_g 0.000373079f
cc_53 N_NET13_20 N_MM5@2_g 0.0331592f
cc_54 N_NET13_18 N_A2_1 0.000583235f
cc_55 N_NET13_20 N_A2_2 0.00079477f
cc_56 N_NET13_5 N_MM5@2_g 0.00104898f
cc_57 N_NET13_18 N_MM5_g 0.0344774f
cc_58 N_NET13_4 N_MM4_g 0.00193786f
cc_59 N_NET13_19 N_A1_1 0.00223976f
cc_60 N_NET13_19 N_MM4@2_g 0.0183757f
cc_61 N_NET13_19 N_MM4_g 0.0497292f
x_PM_AOI22x1_ASAP7_75t_R%Y VSS Y N_MM7@2_d N_MM7_d N_MM6@2_d N_MM6_d N_MM4@2_d
+ N_MM5@2_d N_MM5_d N_MM4_d N_Y_1 N_Y_17 N_Y_2 N_Y_16 N_Y_21 N_Y_20 N_Y_19
+ N_Y_3 N_Y_4 N_Y_5 N_Y_23 N_Y_22 N_Y_18 N_Y_25 PM_AOI22x1_ASAP7_75t_R%Y
cc_62 N_Y_1 N_MM7@2_g 0.00232642f
cc_63 N_Y_17 N_MM3@2_g 0.0345158f
cc_64 N_Y_2 N_B2_9 0.000684459f
cc_65 N_Y_17 N_B2_2 0.000754991f
cc_66 N_Y_16 N_B2_1 0.000810793f
cc_67 N_Y_1 N_B2_7 0.00086092f
cc_68 N_Y_21 N_B2_10 0.00127443f
cc_69 N_Y_2 N_MM3@2_g 0.00161856f
cc_70 N_Y_21 N_B2_8 0.00532459f
cc_71 N_Y_21 N_B2_12 0.00885772f
cc_72 N_Y_16 N_MM7@2_g 0.0355754f
cc_73 N_Y_20 N_MM5@2_g 0.0153111f
cc_74 N_Y_17 N_MM5@2_g 0.000429427f
cc_75 N_Y_19 N_MM5@2_g 0.000433806f
cc_76 N_Y_3 N_A2_1 0.000523175f
cc_77 N_Y_4 N_A2_2 0.000766684f
cc_78 N_Y_3 N_MM5_g 0.000885847f
cc_79 N_Y_4 N_MM5@2_g 0.00102654f
cc_80 N_Y_2 N_A2_7 0.0010507f
cc_81 N_Y_19 N_A2_1 0.00149762f
cc_82 N_Y_2 N_MM5_g 0.00161718f
cc_83 N_Y_21 N_A2_12 0.00166244f
cc_84 N_Y_20 N_A2_2 0.00171191f
cc_85 N_Y_5 N_MM5@2_g 0.00176573f
cc_86 N_Y_23 N_A2_9 0.00425864f
cc_87 N_Y_22 N_A2_11 0.00515014f
cc_88 N_Y_19 N_MM5_g 0.0148888f
cc_89 N_Y_21 N_A2_8 0.00571419f
cc_90 N_Y_21 N_A2_10 0.00847131f
cc_91 N_Y_17 N_MM5_g 0.0524504f
cc_92 N_Y_18 N_MM5@2_g 0.0539874f
cc_93 N_Y_22 N_MM4@2_g 0.000315478f
cc_94 N_Y_3 N_MM4@2_g 0.000351222f
cc_95 N_Y_19 N_MM4@2_g 0.000437719f
cc_96 N_Y_21 N_MM4@2_g 0.000534328f
cc_97 N_Y_4 N_MM4@2_g 0.000799675f
cc_98 N_Y_3 N_MM4_g 0.000957399f
cc_99 N_Y_20 N_A1_1 0.00196272f
cc_100 N_Y_22 N_A1_7 0.00460388f
cc_101 N_Y_19 N_MM4_g 0.0337194f
cc_102 N_Y_20 N_MM4@2_g 0.0351414f
cc_103 N_Y_16 N_NET13_21 0.000196773f
cc_104 N_Y_1 N_NET13_16 0.00020171f
cc_105 N_Y_16 N_NET13_16 0.000219462f
cc_106 N_Y_3 N_NET13_3 0.00443958f
cc_107 N_Y_22 N_NET13_4 0.000571103f
cc_108 N_Y_4 N_NET13_21 0.000577629f
cc_109 N_Y_19 N_NET13_18 0.00171379f
cc_110 N_Y_25 N_NET13_21 0.000632067f
cc_111 N_Y_22 N_NET13_5 0.000683688f
cc_112 N_Y_3 N_NET13_21 0.000697522f
cc_113 N_Y_23 N_NET13_5 0.000706008f
cc_114 N_Y_20 N_NET13_20 0.000739226f
cc_115 N_Y_19 N_NET13_19 0.00111936f
cc_116 N_Y_20 N_NET13_19 0.00112444f
cc_117 N_Y_4 N_NET13_5 0.00249184f
cc_118 N_Y_4 N_NET13_4 0.00274024f
cc_119 N_Y_3 N_NET13_4 0.00305696f
cc_120 N_Y_22 N_NET13_21 0.0177658f
*END of AOI22x1_ASAP7_75t_R.pxi
.ENDS
** Design:	AOI22xp33_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AOI22xp33_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AOI22xp33_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AOI22xp33_ASAP7_75t_R%NET29 VSS 2 3 1
c1 1 VSS 0.000859804f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0540 $X2=0.2160 $Y2=0.0540
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0540 $X2=0.2160 $Y2=0.0540
.ends

.subckt PM_AOI22xp33_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.032333f
.ends

.subckt PM_AOI22xp33_ASAP7_75t_R%NET30 VSS 2 3 1
c1 1 VSS 0.000853524f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0540 $X2=0.1080 $Y2=0.0540
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0540 $X2=0.1080 $Y2=0.0540
.ends

.subckt PM_AOI22xp33_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.00528114f
.ends

.subckt PM_AOI22xp33_ASAP7_75t_R%B2 VSS 6 3 1 4
c1 1 VSS 0.00513295f
c2 3 VSS 0.00792901f
c3 4 VSS 0.00352414f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1207 $X2=0.1890 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1150 $X2=0.1890 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1150 $X2=0.1890 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AOI22xp33_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00485492f
.ends

.subckt PM_AOI22xp33_ASAP7_75t_R%A1 VSS 8 3 1 4
c1 1 VSS 0.00234488f
c2 3 VSS 0.0608826f
c3 4 VSS 0.0145578f
r1 8 7 4.95528 $w=1.3e-08 $l=2.13e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1860 $X2=0.0810 $Y2=0.1647
r2 6 7 6.9374 $w=1.3e-08 $l=2.97e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1647
r3 4 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0980 $X2=0.0810 $Y2=0.1350
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r5 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AOI22xp33_ASAP7_75t_R%A2 VSS 9 3 1 4
c1 1 VSS 0.00397161f
c2 3 VSS 0.034413f
c3 4 VSS 0.00382364f
r1 9 8 2.62338 $w=1.3e-08 $l=1.13e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1860 $X2=0.1350 $Y2=0.1747
r2 7 8 4.83869 $w=1.3e-08 $l=2.07e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1540 $X2=0.1350 $Y2=0.1747
r3 6 7 4.4306 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1540
r4 4 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0980 $X2=0.1350 $Y2=0.1350
r5 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r6 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AOI22xp33_ASAP7_75t_R%B1 VSS 6 3 1 4
c1 1 VSS 0.00411346f
c2 3 VSS 0.0345878f
c3 4 VSS 0.00327539f
r1 7 8 7.28718 $w=1.3e-08 $l=3.13e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1037 $X2=0.2430 $Y2=0.1350
r2 6 7 5.30507 $w=1.3e-08 $l=2.27e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0810 $X2=0.2430 $Y2=0.1037
r3 6 4 1.34084 $w=1.3e-08 $l=5.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0810 $X2=0.2430 $Y2=0.0752
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AOI22xp33_ASAP7_75t_R%Y VSS 26 16 17 36 37 9 1 7 2 10 8 11 13
c1 1 VSS 0.00675683f
c2 2 VSS 0.00293072f
c3 7 VSS 0.00313592f
c4 8 VSS 0.00213618f
c5 9 VSS 0.0140421f
c6 10 VSS 0.000747094f
c7 11 VSS 0.00353708f
c8 12 VSS 0.00348513f
c9 13 VSS 0.00077977f
r1 37 35 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2160 $X2=0.2305 $Y2=0.2160
r2 2 35 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2160 $X2=0.2305 $Y2=0.2160
r3 8 2 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2160 $X2=0.2160 $Y2=0.2160
r4 36 8 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2160 $X2=0.2015 $Y2=0.2160
r5 2 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2160
+ $X2=0.2160 $Y2=0.1980
r6 32 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1980 $X2=0.2295 $Y2=0.1980
r7 30 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1980 $X2=0.2295 $Y2=0.1980
r8 29 30 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2680
+ $Y=0.1980 $X2=0.2430 $Y2=0.1980
r9 10 13 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2860 $Y=0.1980 $X2=0.2970 $Y2=0.1980
r10 10 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2860
+ $Y=0.1980 $X2=0.2680 $Y2=0.1980
r11 13 28 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1980 $X2=0.2970 $Y2=0.1765
r12 27 28 8.68632 $w=1.3e-08 $l=3.73e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1392 $X2=0.2970 $Y2=0.1765
r13 26 27 5.88804 $w=1.3e-08 $l=2.52e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1140 $X2=0.2970 $Y2=0.1392
r14 26 25 5.18847 $w=1.3e-08 $l=2.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1140 $X2=0.2970 $Y2=0.0917
r15 11 12 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0575 $X2=0.2970 $Y2=0.0360
r16 11 25 7.98675 $w=1.3e-08 $l=3.42e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0575 $X2=0.2970 $Y2=0.0917
r17 12 24 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0360 $X2=0.2700 $Y2=0.0360
r18 23 24 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r19 22 23 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2180
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r20 21 22 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2000
+ $Y=0.0360 $X2=0.2180 $Y2=0.0360
r21 20 21 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.2000 $Y2=0.0360
r22 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1755
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r23 18 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r24 9 18 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1505
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r25 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r26 17 15 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0540 $X2=0.1765 $Y2=0.0540
r27 1 15 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.0540 $X2=0.1765 $Y2=0.0540
r28 7 1 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1620 $Y2=0.0540
r29 16 7 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
.ends

.subckt PM_AOI22xp33_ASAP7_75t_R%NET13 VSS 15 32 33 35 1 13 10 2 11 12 3
c1 1 VSS 0.00751659f
c2 2 VSS 0.006028f
c3 3 VSS 0.00534784f
c4 10 VSS 0.00332379f
c5 11 VSS 0.00294951f
c6 12 VSS 0.00237012f
c7 13 VSS 0.0212052f
r1 12 3 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2160 $X2=0.2680 $Y2=0.2160
r2 35 12 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2160 $X2=0.2555 $Y2=0.2160
r3 33 31 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2160 $X2=0.1765 $Y2=0.2160
r4 2 31 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2160 $X2=0.1765 $Y2=0.2160
r5 11 2 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1620 $Y2=0.2160
r6 32 11 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r7 3 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2160
+ $X2=0.2700 $Y2=0.2340
r8 2 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r9 27 28 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2315
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r10 26 27 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2000
+ $Y=0.2340 $X2=0.2315 $Y2=0.2340
r11 25 26 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.2000 $Y2=0.2340
r12 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1755
+ $Y=0.2340 $X2=0.1890 $Y2=0.2340
r13 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r14 22 23 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1505
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r15 21 22 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1460
+ $Y=0.2340 $X2=0.1505 $Y2=0.2340
r16 20 21 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1460 $Y2=0.2340
r17 19 20 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r18 18 19 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.2340 $X2=0.1080 $Y2=0.2340
r19 17 18 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0675
+ $Y=0.2340 $X2=0.0810 $Y2=0.2340
r20 16 17 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2340 $X2=0.0675 $Y2=0.2340
r21 13 16 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r22 1 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0540 $Y2=0.2340
r23 15 14 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r24 10 14 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r25 1 10 1e-05
.ends

.subckt PM_AOI22xp33_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.0319012f
.ends


*
.SUBCKT AOI22xp33_ASAP7_75t_R VSS VDD A1 A2 B2 B1 Y
*
* VSS VSS
* VDD VDD
* A1 A1
* A2 A2
* B2 B2
* B1 B1
* Y Y
*
*

MM8 N_MM8_d N_MM8_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM6 N_MM6_d N_MM6_g N_MM6_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM7 N_MM7_d N_MM7_g N_MM7_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM9 N_MM9_d N_MM9_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2 N_MM2_d N_MM8_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM6_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM7_g N_MM5_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM4 N_MM4_d N_MM9_g N_MM4_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2


*include "AOI22xp33_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AOI22xp33_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AOI22xp33_ASAP7_75t_R%NET29 VSS N_MM7_s N_MM9_d N_NET29_1
+ PM_AOI22xp33_ASAP7_75t_R%NET29
cc_1 N_NET29_1 N_MM7_g 0.012578f
cc_2 N_NET29_1 N_MM9_g 0.0125249f
x_PM_AOI22xp33_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_AOI22xp33_ASAP7_75t_R%noxref_11
cc_3 N_noxref_11_1 N_MM8_g 0.00401251f
x_PM_AOI22xp33_ASAP7_75t_R%NET30 VSS N_MM8_d N_MM6_s N_NET30_1
+ PM_AOI22xp33_ASAP7_75t_R%NET30
cc_4 N_NET30_1 N_MM8_g 0.0125182f
cc_5 N_NET30_1 N_MM6_g 0.0124526f
x_PM_AOI22xp33_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_AOI22xp33_ASAP7_75t_R%noxref_12
cc_6 N_noxref_12_1 N_MM8_g 0.00396006f
cc_7 N_noxref_12_1 N_NET13_10 0.0270924f
cc_8 N_noxref_12_1 N_noxref_11_1 0.00208528f
x_PM_AOI22xp33_ASAP7_75t_R%B2 VSS B2 N_MM7_g N_B2_1 N_B2_4
+ PM_AOI22xp33_ASAP7_75t_R%B2
cc_9 N_B2_1 N_A2_1 0.00166725f
cc_10 N_B2_4 N_A2_4 0.00401951f
cc_11 N_MM7_g N_MM6_g 0.00843545f
x_PM_AOI22xp33_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_AOI22xp33_ASAP7_75t_R%noxref_14
cc_12 N_noxref_14_1 N_MM9_g 0.00366941f
cc_13 N_noxref_14_1 N_NET13_12 0.0270813f
cc_14 N_noxref_14_1 N_Y_8 0.000920265f
cc_15 N_noxref_14_1 N_noxref_13_1 0.00205145f
x_PM_AOI22xp33_ASAP7_75t_R%A1 VSS A1 N_MM8_g N_A1_1 N_A1_4
+ PM_AOI22xp33_ASAP7_75t_R%A1
x_PM_AOI22xp33_ASAP7_75t_R%A2 VSS A2 N_MM6_g N_A2_1 N_A2_4
+ PM_AOI22xp33_ASAP7_75t_R%A2
cc_16 N_A2_1 N_A1_1 0.00161129f
cc_17 N_A2_4 N_A1_4 0.00554806f
cc_18 N_MM6_g N_MM8_g 0.00997462f
x_PM_AOI22xp33_ASAP7_75t_R%B1 VSS B1 N_MM9_g N_B1_1 N_B1_4
+ PM_AOI22xp33_ASAP7_75t_R%B1
cc_19 N_B1_1 N_B2_1 0.00175649f
cc_20 N_B1_4 N_B2_4 0.00368452f
cc_21 N_MM9_g N_MM7_g 0.00978442f
x_PM_AOI22xp33_ASAP7_75t_R%Y VSS Y N_MM6_d N_MM7_d N_MM5_d N_MM4_d N_Y_9 N_Y_1
+ N_Y_7 N_Y_2 N_Y_10 N_Y_8 N_Y_11 N_Y_13 PM_AOI22xp33_ASAP7_75t_R%Y
cc_22 N_Y_9 N_A2_4 0.000561211f
cc_23 N_Y_1 N_MM6_g 0.000966204f
cc_24 N_Y_1 N_A2_4 0.00128575f
cc_25 N_Y_7 N_MM6_g 0.0263781f
cc_26 N_Y_2 N_MM7_g 0.000479248f
cc_27 N_Y_10 N_B2_4 0.000596258f
cc_28 N_Y_8 N_B2_1 0.000634254f
cc_29 N_Y_1 N_MM7_g 0.000946508f
cc_30 N_Y_9 N_B2_4 0.00122761f
cc_31 N_Y_1 N_B2_4 0.00254455f
cc_32 N_Y_8 N_MM7_g 0.0109775f
cc_33 N_Y_7 N_MM7_g 0.0402269f
cc_34 N_Y_11 N_B1_1 0.000555611f
cc_35 N_Y_8 N_B1_1 0.00063387f
cc_36 N_Y_10 N_B1_4 0.00118564f
cc_37 N_Y_9 N_B1_4 0.0012036f
cc_38 N_Y_11 N_B1_4 0.00617745f
cc_39 N_Y_8 N_MM9_g 0.0263413f
cc_40 N_Y_8 N_NET13_12 0.000520211f
cc_41 N_Y_13 N_NET13_13 0.000586418f
cc_42 N_Y_10 N_NET13_3 0.00067674f
cc_43 N_Y_2 N_NET13_13 0.000678327f
cc_44 N_Y_8 N_NET13_11 0.000842661f
cc_45 N_Y_2 N_NET13_3 0.00171401f
cc_46 N_Y_2 N_NET13_2 0.00312627f
cc_47 N_Y_10 N_NET13_13 0.00907101f
x_PM_AOI22xp33_ASAP7_75t_R%NET13 VSS N_MM2_d N_MM3_d N_MM5_s N_MM4_s N_NET13_1
+ N_NET13_13 N_NET13_10 N_NET13_2 N_NET13_11 N_NET13_12 N_NET13_3
+ PM_AOI22xp33_ASAP7_75t_R%NET13
cc_48 N_NET13_1 N_MM8_g 0.000886113f
cc_49 N_NET13_13 N_A1_4 0.00135133f
cc_50 N_NET13_1 N_A1_4 0.00188022f
cc_51 N_NET13_10 N_MM8_g 0.0254499f
cc_52 N_NET13_13 N_A2_4 0.00127026f
cc_53 N_NET13_2 N_A2_4 0.00163646f
cc_54 N_NET13_11 N_MM6_g 0.0258699f
cc_55 N_NET13_2 N_MM7_g 0.000480122f
cc_56 N_NET13_11 N_MM7_g 0.0255831f
cc_57 N_NET13_12 N_MM9_g 0.0259097f
x_PM_AOI22xp33_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_AOI22xp33_ASAP7_75t_R%noxref_13
cc_58 N_noxref_13_1 N_MM9_g 0.00369279f
cc_59 N_noxref_13_1 N_Y_11 0.000937723f
*END of AOI22xp33_ASAP7_75t_R.pxi
.ENDS
** Design:	AOI22xp5_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AOI22xp5_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AOI22xp5_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AOI22xp5_ASAP7_75t_R%NET29 VSS 2 3 1
c1 1 VSS 0.0010082f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2160 $Y2=0.0675
.ends

.subckt PM_AOI22xp5_ASAP7_75t_R%NET30 VSS 2 3 1
c1 1 VSS 0.00100378f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_AOI22xp5_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.00635508f
.ends

.subckt PM_AOI22xp5_ASAP7_75t_R%A1 VSS 15 3 1 6 5 9
c1 1 VSS 0.00425813f
c2 3 VSS 0.0821966f
c3 4 VSS 0.00782594f
c4 5 VSS 0.00310988f
c5 6 VSS 0.0024903f
c6 7 VSS 0.00855568f
c7 8 VSS 0.00156248f
c8 9 VSS 0.00293497f
r1 9 16 5.29071 $w=1.46216e-08 $l=2.78e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1980 $X2=0.0270 $Y2=0.1702
r2 7 14 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0360 $X2=0.0270 $Y2=0.0575
r3 15 16 4.4889 $w=1.3e-08 $l=1.92e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1510 $X2=0.0270 $Y2=0.1702
r4 15 5 0.874462 $w=1.3e-08 $l=3.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1510 $X2=0.0270 $Y2=0.1472
r5 5 8 1.67627 $w=1.66735e-08 $l=1.22e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1472 $X2=0.0270 $Y2=0.1350
r6 4 8 7.44771 $w=1.42162e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0980 $X2=0.0270 $Y2=0.1350
r7 4 14 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0980 $X2=0.0270 $Y2=0.0575
r8 8 13 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1350 $X2=0.0455 $Y2=0.1350
r9 6 11 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.0635
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r10 6 13 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0635
+ $Y=0.1350 $X2=0.0455 $Y2=0.1350
r11 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r12 1 11 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AOI22xp5_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.0419502f
.ends

.subckt PM_AOI22xp5_ASAP7_75t_R%B2 VSS 6 3 1 4
c1 1 VSS 0.00754007f
c2 3 VSS 0.00917647f
c3 4 VSS 0.0046201f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1207 $X2=0.1890 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1150 $X2=0.1890 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1150 $X2=0.1890 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AOI22xp5_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.0418299f
.ends

.subckt PM_AOI22xp5_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00627908f
.ends

.subckt PM_AOI22xp5_ASAP7_75t_R%Y VSS 26 16 17 36 37 9 7 1 10 2 8 11
c1 1 VSS 0.0067481f
c2 2 VSS 0.00291608f
c3 7 VSS 0.00324935f
c4 8 VSS 0.002144f
c5 9 VSS 0.0143886f
c6 10 VSS 0.000656627f
c7 11 VSS 0.00399085f
c8 12 VSS 0.00338888f
c9 13 VSS 0.000784169f
r1 37 35 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r2 2 35 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r4 36 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r5 2 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.1980
r6 32 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1980 $X2=0.2295 $Y2=0.1980
r7 30 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1980 $X2=0.2295 $Y2=0.1980
r8 29 30 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2680
+ $Y=0.1980 $X2=0.2430 $Y2=0.1980
r9 10 13 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2860 $Y=0.1980 $X2=0.2970 $Y2=0.1980
r10 10 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2860
+ $Y=0.1980 $X2=0.2680 $Y2=0.1980
r11 13 28 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1980 $X2=0.2970 $Y2=0.1765
r12 27 28 8.68632 $w=1.3e-08 $l=3.73e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1392 $X2=0.2970 $Y2=0.1765
r13 26 27 5.88804 $w=1.3e-08 $l=2.52e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1140 $X2=0.2970 $Y2=0.1392
r14 26 25 5.18847 $w=1.3e-08 $l=2.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1140 $X2=0.2970 $Y2=0.0917
r15 11 12 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0575 $X2=0.2970 $Y2=0.0360
r16 11 25 7.98675 $w=1.3e-08 $l=3.42e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0575 $X2=0.2970 $Y2=0.0917
r17 12 24 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0360 $X2=0.2700 $Y2=0.0360
r18 23 24 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r19 22 23 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2180
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r20 21 22 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2000
+ $Y=0.0360 $X2=0.2180 $Y2=0.0360
r21 20 21 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.2000 $Y2=0.0360
r22 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1755
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r23 18 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r24 9 18 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1505
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r25 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0675
+ $X2=0.1620 $Y2=0.0360
r26 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r27 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r28 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r29 16 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1475 $Y2=0.0675
.ends

.subckt PM_AOI22xp5_ASAP7_75t_R%B1 VSS 6 3 1 4
c1 1 VSS 0.00716333f
c2 3 VSS 0.0462816f
c3 4 VSS 0.00460909f
r1 7 8 7.28718 $w=1.3e-08 $l=3.13e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1037 $X2=0.2430 $Y2=0.1350
r2 6 7 5.30507 $w=1.3e-08 $l=2.27e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0810 $X2=0.2430 $Y2=0.1037
r3 6 4 1.34084 $w=1.3e-08 $l=5.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0810 $X2=0.2430 $Y2=0.0752
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AOI22xp5_ASAP7_75t_R%A2 VSS 10 3 1 4 5
c1 1 VSS 0.00707005f
c2 3 VSS 0.0457991f
c3 4 VSS 0.00485571f
c4 5 VSS 0.00369177f
r1 5 11 1.20989 $w=1.73902e-08 $l=1.03e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1980 $X2=0.1350 $Y2=0.1877
r2 10 11 0.408082 $w=1.3e-08 $l=1.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1860 $X2=0.1350 $Y2=0.1877
r3 10 9 2.62338 $w=1.3e-08 $l=1.13e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1860 $X2=0.1350 $Y2=0.1747
r4 8 9 4.83869 $w=1.3e-08 $l=2.07e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1540 $X2=0.1350 $Y2=0.1747
r5 4 8 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1540
r6 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r7 1 4 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AOI22xp5_ASAP7_75t_R%NET13 VSS 15 32 33 35 1 10 13 2 11 12 3
c1 1 VSS 0.0078828f
c2 2 VSS 0.00696505f
c3 3 VSS 0.00549502f
c4 10 VSS 0.00371688f
c5 11 VSS 0.00323061f
c6 12 VSS 0.00248765f
c7 13 VSS 0.0201091f
r1 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2680 $Y2=0.2025
r2 35 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r3 33 31 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r4 2 31 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r5 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r6 32 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r7 3 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.2340
r8 2 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r9 27 28 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2315
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r10 26 27 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2000
+ $Y=0.2340 $X2=0.2315 $Y2=0.2340
r11 25 26 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.2000 $Y2=0.2340
r12 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1755
+ $Y=0.2340 $X2=0.1890 $Y2=0.2340
r13 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r14 22 23 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1505
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r15 21 22 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1460
+ $Y=0.2340 $X2=0.1505 $Y2=0.2340
r16 20 21 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1255
+ $Y=0.2340 $X2=0.1460 $Y2=0.2340
r17 19 20 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1010
+ $Y=0.2340 $X2=0.1255 $Y2=0.2340
r18 18 19 5.13017 $w=1.3e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0790
+ $Y=0.2340 $X2=0.1010 $Y2=0.2340
r19 17 18 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0590
+ $Y=0.2340 $X2=0.0790 $Y2=0.2340
r20 16 17 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0500
+ $Y=0.2340 $X2=0.0590 $Y2=0.2340
r21 13 16 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.2340 $X2=0.0500 $Y2=0.2340
r22 1 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0500 $Y2=0.2340
r23 15 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r24 10 14 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r25 1 10 1e-05
.ends


*
.SUBCKT AOI22xp5_ASAP7_75t_R VSS VDD A1 A2 B2 B1 Y
*
* VSS VSS
* VDD VDD
* A1 A1
* A2 A2
* B2 B2
* B1 B1
* Y Y
*
*

MM8 N_MM8_d N_MM8_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM6_g N_MM6_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM7_g N_MM7_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM8_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM6_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM7_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM9_g N_MM4_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AOI22xp5_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AOI22xp5_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AOI22xp5_ASAP7_75t_R%NET29 VSS N_MM7_s N_MM9_d N_NET29_1
+ PM_AOI22xp5_ASAP7_75t_R%NET29
cc_1 N_NET29_1 N_MM7_g 0.0173571f
cc_2 N_NET29_1 N_MM9_g 0.0174354f
x_PM_AOI22xp5_ASAP7_75t_R%NET30 VSS N_MM8_d N_MM6_s N_NET30_1
+ PM_AOI22xp5_ASAP7_75t_R%NET30
cc_3 N_NET30_1 N_MM8_g 0.017193f
cc_4 N_NET30_1 N_MM6_g 0.0173703f
x_PM_AOI22xp5_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_AOI22xp5_ASAP7_75t_R%noxref_12
cc_5 N_noxref_12_1 N_MM8_g 0.00213929f
cc_6 N_noxref_12_1 N_NET13_10 0.0361848f
cc_7 N_noxref_12_1 N_noxref_11_1 0.00176418f
x_PM_AOI22xp5_ASAP7_75t_R%A1 VSS A1 N_MM8_g N_A1_1 N_A1_6 N_A1_5 N_A1_9
+ PM_AOI22xp5_ASAP7_75t_R%A1
x_PM_AOI22xp5_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_AOI22xp5_ASAP7_75t_R%noxref_11
cc_8 N_noxref_11_1 N_MM8_g 0.00224129f
cc_9 N_noxref_11_1 N_NET13_10 0.000475513f
x_PM_AOI22xp5_ASAP7_75t_R%B2 VSS B2 N_MM7_g N_B2_1 N_B2_4
+ PM_AOI22xp5_ASAP7_75t_R%B2
cc_10 N_B2_1 N_A2_1 0.000872931f
cc_11 N_MM7_g N_MM6_g 0.00328339f
cc_12 N_B2_4 N_A2_4 0.00472016f
x_PM_AOI22xp5_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_AOI22xp5_ASAP7_75t_R%noxref_13
cc_13 N_noxref_13_1 N_MM9_g 0.00145093f
cc_14 N_noxref_13_1 N_NET13_12 0.000474279f
cc_15 N_noxref_13_1 N_Y_11 0.00075829f
x_PM_AOI22xp5_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_AOI22xp5_ASAP7_75t_R%noxref_14
cc_16 N_noxref_14_1 N_MM9_g 0.00144005f
cc_17 N_noxref_14_1 N_NET13_12 0.0362227f
cc_18 N_noxref_14_1 N_Y_8 0.000727833f
cc_19 N_noxref_14_1 N_noxref_13_1 0.00177747f
x_PM_AOI22xp5_ASAP7_75t_R%Y VSS Y N_MM6_d N_MM7_d N_MM5_d N_MM4_d N_Y_9 N_Y_7
+ N_Y_1 N_Y_10 N_Y_2 N_Y_8 N_Y_11 PM_AOI22xp5_ASAP7_75t_R%Y
cc_20 N_Y_9 N_A2_4 0.000604027f
cc_21 N_Y_7 N_A2_1 0.000687241f
cc_22 N_Y_1 N_A2_4 0.00141422f
cc_23 N_Y_1 N_MM6_g 0.00156228f
cc_24 N_Y_7 N_MM6_g 0.0354655f
cc_25 N_Y_7 N_B2_1 0.000502825f
cc_26 N_Y_10 N_B2_4 0.000548857f
cc_27 N_Y_2 N_MM7_g 0.000880385f
cc_28 N_Y_9 N_B2_4 0.00116827f
cc_29 N_Y_1 N_MM7_g 0.00149861f
cc_30 N_Y_8 N_B2_1 0.00154969f
cc_31 N_Y_1 N_B2_4 0.00248886f
cc_32 N_Y_8 N_MM7_g 0.0149884f
cc_33 N_Y_7 N_MM7_g 0.0541101f
cc_34 N_Y_8 N_B1_1 0.00138088f
cc_35 N_Y_2 N_MM9_g 0.000873117f
cc_36 N_Y_10 N_B1_4 0.00106037f
cc_37 N_Y_9 N_B1_4 0.00122063f
cc_38 N_Y_11 N_B1_4 0.00616006f
cc_39 N_Y_8 N_MM9_g 0.0349486f
cc_40 N_Y_10 N_NET13_3 0.000664902f
cc_41 N_Y_8 N_NET13_12 0.00179946f
cc_42 N_Y_11 N_NET13_3 0.00072226f
cc_43 N_Y_2 N_NET13_13 0.000768393f
cc_44 N_Y_2 N_NET13_2 0.00137321f
cc_45 N_Y_2 N_NET13_3 0.0051936f
cc_46 N_Y_10 N_NET13_13 0.00936513f
x_PM_AOI22xp5_ASAP7_75t_R%B1 VSS B1 N_MM9_g N_B1_1 N_B1_4
+ PM_AOI22xp5_ASAP7_75t_R%B1
cc_47 N_B1_1 N_B2_1 0.00114442f
cc_48 N_B1_4 N_B2_4 0.00324761f
cc_49 N_MM9_g N_MM7_g 0.00580973f
x_PM_AOI22xp5_ASAP7_75t_R%A2 VSS A2 N_MM6_g N_A2_1 N_A2_4 N_A2_5
+ PM_AOI22xp5_ASAP7_75t_R%A2
cc_50 N_A2_1 N_A1_1 0.00173896f
cc_51 N_A2_4 N_A1_6 0.00289495f
cc_52 N_MM6_g N_MM8_g 0.00665653f
x_PM_AOI22xp5_ASAP7_75t_R%NET13 VSS N_MM2_d N_MM3_d N_MM5_s N_MM4_s N_NET13_1
+ N_NET13_10 N_NET13_13 N_NET13_2 N_NET13_11 N_NET13_12 N_NET13_3
+ PM_AOI22xp5_ASAP7_75t_R%NET13
cc_53 N_NET13_1 N_A1_5 0.000517358f
cc_54 N_NET13_10 N_A1_1 0.000788274f
cc_55 N_NET13_1 N_MM8_g 0.00197139f
cc_56 N_NET13_13 N_A1_9 0.00332861f
cc_57 N_NET13_10 N_MM8_g 0.0351083f
cc_58 N_NET13_2 N_MM6_g 0.00194253f
cc_59 N_NET13_11 N_A2_1 0.000817616f
cc_60 N_NET13_13 N_A2_5 0.00482643f
cc_61 N_NET13_11 N_MM6_g 0.034179f
cc_62 N_NET13_11 N_B2_1 0.000735789f
cc_63 N_NET13_2 N_MM7_g 0.000940784f
cc_64 N_NET13_11 N_MM7_g 0.0345435f
cc_65 N_NET13_12 N_B1_1 0.000646493f
cc_66 N_NET13_3 N_MM9_g 0.00101756f
cc_67 N_NET13_12 N_MM9_g 0.0344495f
*END of AOI22xp5_ASAP7_75t_R.pxi
.ENDS
** Design:	AOI311xp33_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AOI311xp33_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AOI311xp33_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AOI311xp33_ASAP7_75t_R%NET30 VSS 2 3 1
c1 1 VSS 0.00093792f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_AOI311xp33_ASAP7_75t_R%NET020 VSS 2 3 1
c1 1 VSS 0.000965077f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2700 $Y2=0.2025
.ends

.subckt PM_AOI311xp33_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.0424761f
.ends

.subckt PM_AOI311xp33_ASAP7_75t_R%NET29 VSS 2 3 1
c1 1 VSS 0.000952335f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_AOI311xp33_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.0424937f
.ends

.subckt PM_AOI311xp33_ASAP7_75t_R%NET23 VSS 12 13 24 27 7 1 9 2 8
c1 1 VSS 0.00953528f
c2 2 VSS 0.00841289f
c3 7 VSS 0.00450417f
c4 8 VSS 0.00424661f
c5 9 VSS 0.014344f
r1 27 26 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r2 25 26 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2260 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r3 2 25 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2140 $Y=0.2025 $X2=0.2260 $Y2=0.2025
r4 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2140 $Y2=0.2025
r5 24 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r6 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.2340
r7 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2025
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r8 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.2025 $Y2=0.2340
r9 18 19 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1890 $Y2=0.2340
r10 17 18 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r11 16 17 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1215
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r12 15 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.1215 $Y2=0.2340
r13 14 15 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0970
+ $Y=0.2340 $X2=0.1080 $Y2=0.2340
r14 9 14 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.2340 $X2=0.0970 $Y2=0.2340
r15 1 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.2340
r16 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r17 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r18 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r19 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
.ends

.subckt PM_AOI311xp33_ASAP7_75t_R%A3 VSS 9 3 1 6
c1 1 VSS 0.00482701f
c2 3 VSS 0.0821253f
c3 4 VSS 0.011862f
c4 5 VSS 0.0112514f
c5 6 VSS 0.00302946f
c6 7 VSS 0.00182756f
r1 5 7 7.44771 $w=1.42162e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1720 $X2=0.0270 $Y2=0.1350
r2 4 7 11.6451 $w=1.38182e-08 $l=5.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0800 $X2=0.0270 $Y2=0.1350
r3 9 6 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0540 $Y2=0.1350
r4 6 7 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.1350 $X2=0.0270 $Y2=0.1350
r5 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r6 9 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AOI311xp33_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00447805f
.ends

.subckt PM_AOI311xp33_ASAP7_75t_R%C VSS 6 3 1 4
c1 1 VSS 0.00516398f
c2 3 VSS 0.0349486f
c3 4 VSS 0.00484079f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.0980
r2 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_AOI311xp33_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.0048036f
.ends

.subckt PM_AOI311xp33_ASAP7_75t_R%A1 VSS 6 3 1 4
c1 1 VSS 0.00827397f
c2 3 VSS 0.046237f
c3 4 VSS 0.00567437f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.0980
r2 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AOI311xp33_ASAP7_75t_R%A2 VSS 4 3 1
c1 1 VSS 0.00713158f
c2 3 VSS 0.0467877f
c3 4 VSS 0.00909351f
r1 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r2 4 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AOI311xp33_ASAP7_75t_R%B VSS 6 3 1 4
c1 1 VSS 0.00583537f
c2 3 VSS 0.0350291f
c3 4 VSS 0.0047555f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.0980
r2 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AOI311xp33_ASAP7_75t_R%Y VSS 31 21 22 42 47 1 10 11 15 14 3 2 12 16
c1 1 VSS 0.00775872f
c2 2 VSS 0.00682019f
c3 3 VSS 0.00599651f
c4 10 VSS 0.00320827f
c5 11 VSS 0.000386194f
c6 12 VSS 0.00310923f
c7 13 VSS 5.05396e-20
c8 14 VSS 0.0027416f
c9 15 VSS 0.0135278f
c10 16 VSS 0.00292851f
c11 17 VSS 0.00602344f
c12 18 VSS 0.0028176f
r1 14 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3220 $Y2=0.2025
r2 47 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r3 3 44 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.2340
r4 44 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.2340 $X2=0.3375 $Y2=0.2340
r5 17 40 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.2340 $X2=0.3510 $Y2=0.2125
r6 17 45 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.2340 $X2=0.3375 $Y2=0.2340
r7 12 2 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0540 $X2=0.3220 $Y2=0.0540
r8 42 12 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0540 $X2=0.3095 $Y2=0.0540
r9 39 40 18.0722 $w=1.3e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.2125
r10 16 18 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.0575 $X2=0.3510 $Y2=0.0360
r11 16 39 18.0722 $w=1.3e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0575 $X2=0.3510 $Y2=0.1350
r12 2 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0540
+ $X2=0.3240 $Y2=0.0360
r13 18 38 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.0360 $X2=0.3375 $Y2=0.0360
r14 37 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.0360 $X2=0.3375 $Y2=0.0360
r15 36 37 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3125
+ $Y=0.0360 $X2=0.3240 $Y2=0.0360
r16 35 36 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3080
+ $Y=0.0360 $X2=0.3125 $Y2=0.0360
r17 34 35 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.3080 $Y2=0.0360
r18 33 34 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.2970 $Y2=0.0360
r19 32 33 4.6055 $w=1.3e-08 $l=1.98e-08 $layer=M1 $thickness=3.6e-08 $X=0.2502
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r20 31 32 0.524677 $w=1.3e-08 $l=2.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.2480
+ $Y=0.0360 $X2=0.2502 $Y2=0.0360
r21 31 30 1.69063 $w=1.3e-08 $l=7.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.2480
+ $Y=0.0360 $X2=0.2407 $Y2=0.0360
r22 29 30 2.62338 $w=1.3e-08 $l=1.12e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.0360 $X2=0.2407 $Y2=0.0360
r23 28 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.2295 $Y2=0.0360
r24 15 28 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2025
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r25 11 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0945 $X2=0.2140 $Y2=0.0945
r26 1 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0540
+ $X2=0.2160 $Y2=0.0360
r27 24 25 0.264706 $w=1.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2260 $Y=0.0725 $X2=0.2305 $Y2=0.0725
r28 1 24 0.705882 $w=1.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2140 $Y=0.0725 $X2=0.2260 $Y2=0.0725
r29 13 1 0.735294 $w=1.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0725 $X2=0.2140 $Y2=0.0725
r30 22 20 0.0675676 $w=3.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0455 $X2=0.2305 $Y2=0.0455
r31 1 20 0.391892 $w=3.7e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.0455 $X2=0.2305 $Y2=0.0455
r32 1 25 0.471383 $w=3.35517e-08 $l=3.06472e-08 $layer=N_src_drn
+ $thickness=1e-09 $X=0.2160 $Y=0.0455 $X2=0.2305 $Y2=0.0725
r33 10 1 0.391892 $w=3.7e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0455 $X2=0.2160 $Y2=0.0455
r34 21 10 0.0675676 $w=3.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0455 $X2=0.2015 $Y2=0.0455
.ends


*
.SUBCKT AOI311xp33_ASAP7_75t_R VSS VDD A3 A2 A1 B C Y
*
* VSS VSS
* VDD VDD
* A3 A3
* A2 A2
* A1 A1
* B B
* C C
* Y Y
*
*

MM4 N_MM4_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g N_MM3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM0 N_MM0_d N_MM0_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM10 N_MM10_d N_MM4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM5_g N_MM9_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM0_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AOI311xp33_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AOI311xp33_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AOI311xp33_ASAP7_75t_R%NET30 VSS N_MM3_d N_MM2_s N_NET30_1
+ PM_AOI311xp33_ASAP7_75t_R%NET30
cc_1 N_NET30_1 N_MM3_g 0.0172888f
cc_2 N_NET30_1 N_MM2_g 0.0171479f
x_PM_AOI311xp33_ASAP7_75t_R%NET020 VSS N_MM9_d N_MM1_s N_NET020_1
+ PM_AOI311xp33_ASAP7_75t_R%NET020
cc_3 N_NET020_1 N_MM5_g 0.0173419f
cc_4 N_NET020_1 N_MM0_g 0.0172318f
x_PM_AOI311xp33_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_AOI311xp33_ASAP7_75t_R%noxref_13
cc_5 N_noxref_13_1 N_MM4_g 0.00222235f
x_PM_AOI311xp33_ASAP7_75t_R%NET29 VSS N_MM4_d N_MM3_s N_NET29_1
+ PM_AOI311xp33_ASAP7_75t_R%NET29
cc_6 N_NET29_1 N_MM4_g 0.0173459f
cc_7 N_NET29_1 N_MM3_g 0.017271f
x_PM_AOI311xp33_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_AOI311xp33_ASAP7_75t_R%noxref_14
cc_8 N_noxref_14_1 N_MM4_g 0.0022148f
cc_9 N_noxref_14_1 N_noxref_13_1 0.00177211f
x_PM_AOI311xp33_ASAP7_75t_R%NET23 VSS N_MM10_d N_MM7_d N_MM6_d N_MM9_s
+ N_NET23_7 N_NET23_1 N_NET23_9 N_NET23_2 N_NET23_8
+ PM_AOI311xp33_ASAP7_75t_R%NET23
cc_10 N_NET23_7 N_A3_1 0.000665015f
cc_11 N_NET23_1 N_MM4_g 0.00101184f
cc_12 N_NET23_7 N_MM4_g 0.034486f
cc_13 N_NET23_7 N_A2_1 0.000753369f
cc_14 N_NET23_9 N_A2 0.00114235f
cc_15 N_NET23_1 N_MM3_g 0.00119856f
cc_16 N_NET23_1 N_A2 0.00173422f
cc_17 N_NET23_7 N_MM3_g 0.0335183f
cc_18 N_NET23_9 N_A1_4 0.00109822f
cc_19 N_NET23_2 N_MM2_g 0.00114733f
cc_20 N_NET23_2 N_A1_4 0.00170675f
cc_21 N_NET23_8 N_MM2_g 0.0342563f
cc_22 N_NET23_8 N_B_1 0.000687941f
cc_23 N_NET23_2 N_B_4 0.00123113f
cc_24 N_NET23_2 N_MM5_g 0.00149283f
cc_25 N_NET23_8 N_MM5_g 0.0345334f
x_PM_AOI311xp33_ASAP7_75t_R%A3 VSS A3 N_MM4_g N_A3_1 N_A3_6
+ PM_AOI311xp33_ASAP7_75t_R%A3
x_PM_AOI311xp33_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_AOI311xp33_ASAP7_75t_R%noxref_15
cc_26 N_noxref_15_1 N_MM0_g 0.00350218f
cc_27 N_noxref_15_1 N_Y_12 0.0287209f
x_PM_AOI311xp33_ASAP7_75t_R%C VSS C N_MM0_g N_C_1 N_C_4
+ PM_AOI311xp33_ASAP7_75t_R%C
cc_28 N_C_1 N_B_1 0.00157883f
cc_29 N_C_4 N_B_4 0.00501846f
cc_30 N_MM0_g N_MM5_g 0.00819212f
x_PM_AOI311xp33_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_AOI311xp33_ASAP7_75t_R%noxref_16
cc_31 N_noxref_16_1 N_MM0_g 0.00160899f
cc_32 N_noxref_16_1 N_Y_14 0.0381706f
cc_33 N_noxref_16_1 N_noxref_15_1 0.00190215f
x_PM_AOI311xp33_ASAP7_75t_R%A1 VSS A1 N_MM2_g N_A1_1 N_A1_4
+ PM_AOI311xp33_ASAP7_75t_R%A1
cc_34 N_A1_1 N_A2_1 0.00125612f
cc_35 N_MM2_g N_MM3_g 0.00519176f
cc_36 N_A1_4 N_A2 0.00638661f
x_PM_AOI311xp33_ASAP7_75t_R%A2 VSS A2 N_MM3_g N_A2_1
+ PM_AOI311xp33_ASAP7_75t_R%A2
cc_37 N_A2_1 N_MM4_g 0.000622825f
cc_38 N_A2_1 N_A3_1 0.00134305f
cc_39 N_A2 N_A3_6 0.00321176f
cc_40 N_MM3_g N_MM4_g 0.00635052f
x_PM_AOI311xp33_ASAP7_75t_R%B VSS B N_MM5_g N_B_1 N_B_4
+ PM_AOI311xp33_ASAP7_75t_R%B
cc_41 N_B_1 N_A1_4 0.000864619f
cc_42 N_MM5_g N_MM2_g 0.00329257f
cc_43 N_B_4 N_A1_4 0.00555965f
x_PM_AOI311xp33_ASAP7_75t_R%Y VSS Y N_MM2_d N_MM5_d N_MM0_d N_MM1_d N_Y_1
+ N_Y_10 N_Y_11 N_Y_15 N_Y_14 N_Y_3 N_Y_2 N_Y_12 N_Y_16
+ PM_AOI311xp33_ASAP7_75t_R%Y
cc_44 N_Y_1 N_A2 0.00171847f
cc_45 N_Y_10 N_A1_1 0.000654597f
cc_46 N_Y_1 N_A1_4 0.00132759f
cc_47 N_Y_1 N_MM2_g 0.00154778f
cc_48 N_Y_10 N_MM2_g 0.00990792f
cc_49 N_Y_11 N_MM2_g 0.0257406f
cc_50 N_Y_10 N_B_1 0.00121297f
cc_51 N_Y_15 N_B_4 0.00112444f
cc_52 N_Y_1 N_MM5_g 0.00130808f
cc_53 N_Y_1 N_B_4 0.0019727f
cc_54 N_Y_11 N_MM5_g 0.00526638f
cc_55 N_Y_10 N_MM5_g 0.0309028f
cc_56 N_Y_14 N_C_4 0.000564919f
cc_57 N_Y_3 N_C_1 0.000678966f
cc_58 N_Y_2 N_MM0_g 0.00075325f
cc_59 N_Y_15 N_C_4 0.00110578f
cc_60 N_Y_14 N_C_1 0.00129075f
cc_61 N_Y_3 N_MM0_g 0.00172992f
cc_62 N_Y_12 N_MM0_g 0.0108902f
cc_63 N_Y_16 N_C_4 0.00796355f
cc_64 N_Y_14 N_MM0_g 0.0501254f
*END of AOI311xp33_ASAP7_75t_R.pxi
.ENDS
** Design:	AOI31xp33_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AOI31xp33_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AOI31xp33_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AOI31xp33_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.0425245f
.ends

.subckt PM_AOI31xp33_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.0327766f
.ends

.subckt PM_AOI31xp33_ASAP7_75t_R%NET30 VSS 2 3 1
c1 1 VSS 0.000910649f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_AOI31xp33_ASAP7_75t_R%A3 VSS 8 3 1 4
c1 1 VSS 0.00419703f
c2 3 VSS 0.0715354f
c3 4 VSS 0.0165401f
r1 8 4 12.7088 $w=1.3e-08 $l=5.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1340 $X2=0.0810 $Y2=0.0795
r2 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1340
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AOI31xp33_ASAP7_75t_R%NET29 VSS 2 3 1
c1 1 VSS 0.000883511f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_AOI31xp33_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00468189f
.ends

.subckt PM_AOI31xp33_ASAP7_75t_R%NET23 VSS 12 13 24 27 1 7 9 2 8
c1 1 VSS 0.00840038f
c2 2 VSS 0.00619775f
c3 7 VSS 0.0038885f
c4 8 VSS 0.00299872f
c5 9 VSS 0.0137367f
r1 27 26 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2160 $X2=0.2305 $Y2=0.2160
r2 25 26 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2260 $Y=0.2160 $X2=0.2305 $Y2=0.2160
r3 2 25 0.222222 $w=5.4e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2140 $Y=0.2160 $X2=0.2260 $Y2=0.2160
r4 8 2 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2160 $X2=0.2140 $Y2=0.2160
r5 24 8 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2160 $X2=0.2015 $Y2=0.2160
r6 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2160
+ $X2=0.2160 $Y2=0.2340
r7 20 21 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2040
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r8 19 20 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1995
+ $Y=0.2340 $X2=0.2040 $Y2=0.2340
r9 18 19 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.1995 $Y2=0.2340
r10 17 18 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1890 $Y2=0.2340
r11 16 17 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r12 15 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1215
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r13 14 15 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.1215 $Y2=0.2340
r14 9 14 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0960
+ $Y=0.2340 $X2=0.1080 $Y2=0.2340
r15 1 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2160
+ $X2=0.1080 $Y2=0.2340
r16 13 11 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2160 $X2=0.1225 $Y2=0.2160
r17 1 11 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2160 $X2=0.1225 $Y2=0.2160
r18 7 1 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2160 $X2=0.1080 $Y2=0.2160
r19 12 7 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2160 $X2=0.0935 $Y2=0.2160
.ends

.subckt PM_AOI31xp33_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.0316723f
.ends

.subckt PM_AOI31xp33_ASAP7_75t_R%B VSS 8 3 1 4
c1 1 VSS 0.00540012f
c2 3 VSS 0.0340814f
c3 4 VSS 0.00380845f
r1 8 4 8.51143 $w=1.3e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1340 $X2=0.2430 $Y2=0.0975
r2 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1340
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AOI31xp33_ASAP7_75t_R%A2 VSS 8 3 1 4
c1 1 VSS 0.00478648f
c2 3 VSS 0.0356317f
c3 4 VSS 0.00734706f
r1 8 4 8.51143 $w=1.3e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1340 $X2=0.1350 $Y2=0.0975
r2 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1340
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AOI31xp33_ASAP7_75t_R%A1 VSS 8 3 1 4
c1 1 VSS 0.00537133f
c2 3 VSS 0.0349032f
c3 4 VSS 0.00461141f
r1 8 4 8.51143 $w=1.3e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1340 $X2=0.1890 $Y2=0.0975
r2 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1340
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AOI31xp33_ASAP7_75t_R%Y VSS 31 17 18 38 1 11 7 8 2 13 10 12
c1 1 VSS 0.00785937f
c2 2 VSS 0.00409648f
c3 7 VSS 0.00306177f
c4 8 VSS 0.000371616f
c5 9 VSS 5.43015e-20
c6 10 VSS 0.00230785f
c7 11 VSS 0.00907856f
c8 12 VSS 0.00350843f
c9 13 VSS 0.0019612f
c10 14 VSS 0.00342829f
r1 10 2 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2160 $X2=0.2680 $Y2=0.2160
r2 38 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2160 $X2=0.2555 $Y2=0.2160
r3 2 35 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2160
+ $X2=0.2700 $Y2=0.1980
r4 35 36 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1980 $X2=0.2835 $Y2=0.1980
r5 13 33 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1980 $X2=0.2970 $Y2=0.1765
r6 13 36 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1980 $X2=0.2835 $Y2=0.1980
r7 32 33 9.0361 $w=1.3e-08 $l=3.88e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1377 $X2=0.2970 $Y2=0.1765
r8 31 32 6.23783 $w=1.3e-08 $l=2.67e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1110 $X2=0.2970 $Y2=0.1377
r9 31 30 4.83869 $w=1.3e-08 $l=2.08e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1110 $X2=0.2970 $Y2=0.0902
r10 12 14 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0575 $X2=0.2970 $Y2=0.0360
r11 12 30 7.63696 $w=1.3e-08 $l=3.27e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0575 $X2=0.2970 $Y2=0.0902
r12 14 29 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.2720 $Y2=0.0360
r13 28 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2540
+ $Y=0.0360 $X2=0.2720 $Y2=0.0360
r14 27 28 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2540 $Y2=0.0360
r15 26 27 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2320
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r16 25 26 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2275
+ $Y=0.0360 $X2=0.2320 $Y2=0.0360
r17 24 25 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.2275 $Y2=0.0360
r18 11 24 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2040
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r19 8 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0945 $X2=0.2140 $Y2=0.0945
r20 1 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0540
+ $X2=0.2160 $Y2=0.0360
r21 20 21 0.264706 $w=1.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2260 $Y=0.0725 $X2=0.2305 $Y2=0.0725
r22 1 20 0.705882 $w=1.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2140 $Y=0.0725 $X2=0.2260 $Y2=0.0725
r23 9 1 0.735294 $w=1.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0725 $X2=0.2140 $Y2=0.0725
r24 18 16 0.0675676 $w=3.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0455 $X2=0.2305 $Y2=0.0455
r25 1 16 0.391892 $w=3.7e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.0455 $X2=0.2305 $Y2=0.0455
r26 1 21 0.471383 $w=3.35517e-08 $l=3.06472e-08 $layer=N_src_drn
+ $thickness=1e-09 $X=0.2160 $Y=0.0455 $X2=0.2305 $Y2=0.0725
r27 7 1 0.391892 $w=3.7e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0455 $X2=0.2160 $Y2=0.0455
r28 17 7 0.0675676 $w=3.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0455 $X2=0.2015 $Y2=0.0455
.ends


*
.SUBCKT AOI31xp33_ASAP7_75t_R VSS VDD A3 A2 A1 B Y
*
* VSS VSS
* VDD VDD
* A3 A3
* A2 A2
* A1 A1
* B B
* Y Y
*
*

MM4 N_MM4_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g N_MM3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM10 N_MM10_d N_MM4_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM7 N_MM7_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM6 N_MM6_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM9 N_MM9_d N_MM5_g N_MM9_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2


*include "AOI31xp33_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AOI31xp33_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AOI31xp33_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_AOI31xp33_ASAP7_75t_R%noxref_11
cc_1 N_noxref_11_1 N_MM4_g 0.00185041f
x_PM_AOI31xp33_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_AOI31xp33_ASAP7_75t_R%noxref_12
cc_2 N_noxref_12_1 N_MM4_g 0.0037631f
cc_3 N_noxref_12_1 N_noxref_11_1 0.00192502f
x_PM_AOI31xp33_ASAP7_75t_R%NET30 VSS N_MM3_d N_MM2_s N_NET30_1
+ PM_AOI31xp33_ASAP7_75t_R%NET30
cc_4 N_NET30_1 N_MM3_g 0.0174704f
cc_5 N_NET30_1 N_MM2_g 0.017283f
x_PM_AOI31xp33_ASAP7_75t_R%A3 VSS A3 N_MM4_g N_A3_1 N_A3_4
+ PM_AOI31xp33_ASAP7_75t_R%A3
x_PM_AOI31xp33_ASAP7_75t_R%NET29 VSS N_MM4_d N_MM3_s N_NET29_1
+ PM_AOI31xp33_ASAP7_75t_R%NET29
cc_6 N_NET29_1 N_MM4_g 0.0172564f
cc_7 N_NET29_1 N_MM3_g 0.0172562f
x_PM_AOI31xp33_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_AOI31xp33_ASAP7_75t_R%noxref_14
cc_8 N_noxref_14_1 N_MM5_g 0.0036564f
cc_9 N_noxref_14_1 N_Y_10 0.0281887f
cc_10 N_noxref_14_1 N_noxref_13_1 0.00205195f
x_PM_AOI31xp33_ASAP7_75t_R%NET23 VSS N_MM10_d N_MM7_d N_MM6_d N_MM9_s N_NET23_1
+ N_NET23_7 N_NET23_9 N_NET23_2 N_NET23_8 PM_AOI31xp33_ASAP7_75t_R%NET23
cc_11 N_NET23_1 N_MM4_g 0.000685291f
cc_12 N_NET23_1 N_A3_4 0.00109951f
cc_13 N_NET23_7 N_MM4_g 0.0253182f
cc_14 N_NET23_1 N_MM3_g 0.000652601f
cc_15 N_NET23_9 N_A2_4 0.00116241f
cc_16 N_NET23_1 N_A2_4 0.00144377f
cc_17 N_NET23_7 N_MM3_g 0.0247151f
cc_18 N_NET23_2 N_MM2_g 0.000708047f
cc_19 N_NET23_9 N_A1_4 0.00123664f
cc_20 N_NET23_2 N_A1_4 0.0016387f
cc_21 N_NET23_8 N_MM2_g 0.024868f
cc_22 N_NET23_2 N_MM5_g 0.000542459f
cc_23 N_NET23_8 N_MM5_g 0.0248383f
x_PM_AOI31xp33_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_AOI31xp33_ASAP7_75t_R%noxref_13
cc_24 N_noxref_13_1 N_MM5_g 0.00364919f
cc_25 N_noxref_13_1 N_Y_8 0.00120429f
x_PM_AOI31xp33_ASAP7_75t_R%B VSS B N_MM5_g N_B_1 N_B_4
+ PM_AOI31xp33_ASAP7_75t_R%B
cc_26 N_B_1 N_A1_1 0.00112513f
cc_27 N_B_4 N_A1_4 0.00401883f
cc_28 N_MM5_g N_MM2_g 0.0063373f
x_PM_AOI31xp33_ASAP7_75t_R%A2 VSS A2 N_MM3_g N_A2_1 N_A2_4
+ PM_AOI31xp33_ASAP7_75t_R%A2
cc_29 N_A2_1 N_A3_1 0.00174409f
cc_30 N_A2_4 N_A3_4 0.00654519f
cc_31 N_MM3_g N_MM4_g 0.00839277f
x_PM_AOI31xp33_ASAP7_75t_R%A1 VSS A1 N_MM2_g N_A1_1 N_A1_4
+ PM_AOI31xp33_ASAP7_75t_R%A1
cc_32 N_A1_1 N_A2_1 0.00161868f
cc_33 N_A1_4 N_A2_4 0.00544763f
cc_34 N_MM2_g N_MM3_g 0.00825434f
x_PM_AOI31xp33_ASAP7_75t_R%Y VSS Y N_MM2_d N_MM5_d N_MM9_d N_Y_1 N_Y_11 N_Y_7
+ N_Y_8 N_Y_2 N_Y_13 N_Y_10 N_Y_12 PM_AOI31xp33_ASAP7_75t_R%Y
cc_35 N_Y_1 N_MM3_g 0.000345041f
cc_36 N_Y_1 N_A2_4 0.00138179f
cc_37 N_Y_11 N_A1_4 0.000543147f
cc_38 N_Y_7 N_A1_1 0.000683282f
cc_39 N_Y_1 N_MM2_g 0.00158309f
cc_40 N_Y_1 N_A1_4 0.00161217f
cc_41 N_Y_7 N_MM2_g 0.0099525f
cc_42 N_Y_8 N_MM2_g 0.0258321f
cc_43 N_Y_2 N_MM5_g 0.000480379f
cc_44 N_Y_13 N_B_4 0.000576022f
cc_45 N_Y_1 N_B_1 0.00077375f
cc_46 N_Y_11 N_B_4 0.00101763f
cc_47 N_Y_7 N_B_1 0.00124012f
cc_48 N_Y_1 N_MM5_g 0.00135293f
cc_49 N_Y_10 N_MM5_g 0.0108773f
cc_50 N_Y_8 N_MM5_g 0.00527887f
cc_51 N_Y_12 N_B_4 0.0064157f
cc_52 N_Y_7 N_MM5_g 0.044462f
cc_53 N_Y_10 N_NET23_8 0.000426296f
cc_54 N_Y_13 N_NET23_9 0.00111536f
cc_55 N_Y_2 N_NET23_2 0.00318461f
*END of AOI31xp33_ASAP7_75t_R.pxi
.ENDS
** Design:	AOI31xp67_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AOI31xp67_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AOI31xp67_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AOI31xp67_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.00647274f
.ends

.subckt PM_AOI31xp67_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00694689f
.ends

.subckt PM_AOI31xp67_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.0417377f
.ends

.subckt PM_AOI31xp67_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.0419599f
.ends

.subckt PM_AOI31xp67_ASAP7_75t_R%A3 VSS 21 3 4 7 1 10
c1 1 VSS 0.00880954f
c2 3 VSS 0.0804547f
c3 4 VSS 0.0803338f
c4 5 VSS 0.0114433f
c5 6 VSS 0.00541365f
c6 7 VSS 0.00323478f
c7 8 VSS 0.00995033f
c8 9 VSS 0.00283343f
c9 10 VSS 0.00501279f
r1 8 27 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0360 $X2=0.0270 $Y2=0.0540
r2 6 9 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1665 $X2=0.0270 $Y2=0.1350
r3 6 10 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1665 $X2=0.0270 $Y2=0.1980
r4 26 27 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0720 $X2=0.0270 $Y2=0.0540
r5 5 9 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1035 $X2=0.0270 $Y2=0.1350
r6 5 26 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1035 $X2=0.0270 $Y2=0.0720
r7 9 23 3.60008 $w=1.51951e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1350 $X2=0.0475 $Y2=0.1350
r8 4 19 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r9 21 7 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0655 $Y2=0.1350
r10 7 23 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0655
+ $Y=0.1350 $X2=0.0475 $Y2=0.1350
r11 17 19 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1350 $X2=0.1350 $Y2=0.1350
r12 16 17 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1350 $X2=0.1225 $Y2=0.1350
r13 15 16 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1350 $X2=0.1080 $Y2=0.1350
r14 13 15 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0905 $Y=0.1350 $X2=0.0935 $Y2=0.1350
r15 12 13 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0905 $Y2=0.1350
r16 21 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
r17 1 12 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r18 1 14 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1350 $X2=0.0705 $Y2=0.1350
r19 3 12 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0810 $Y2=0.1350
r20 3 14 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.0810 $Y=0.1350 $X2=0.0705 $Y2=0.1350
r21 3 15 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1350
.ends

.subckt PM_AOI31xp67_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.00413667f
.ends

.subckt PM_AOI31xp67_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.00416313f
.ends

.subckt PM_AOI31xp67_ASAP7_75t_R%B VSS 21 3 4 8 5 6 10 1 9 7
c1 1 VSS 0.00830766f
c2 3 VSS 0.0448559f
c3 4 VSS 0.00821447f
c4 5 VSS 0.00333801f
c5 6 VSS 0.00316976f
c6 7 VSS 0.00314936f
c7 8 VSS 0.00353669f
c8 9 VSS 0.00376666f
c9 10 VSS 0.00253154f
r1 6 10 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1665 $X2=0.1350 $Y2=0.1350
r2 6 9 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1665 $X2=0.1350 $Y2=0.1980
r3 5 10 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1035 $X2=0.1350 $Y2=0.1350
r4 5 8 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1035 $X2=0.1350 $Y2=0.0720
r5 21 7 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1620 $Y2=0.1350
r6 7 10 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1620 $Y=0.1350 $X2=0.1350 $Y2=0.1350
r7 3 16 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r8 16 17 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1985 $Y2=0.1350
r9 21 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
r10 13 17 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.2015 $Y=0.1350 $X2=0.1985 $Y2=0.1350
r11 12 13 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2160 $Y=0.1350 $X2=0.2015 $Y2=0.1350
r12 11 12 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2305 $Y=0.1350 $X2=0.2160 $Y2=0.1350
r13 4 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r14 1 11 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2305 $Y2=0.1350
r15 1 19 2.90696 $w=2.1681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2535 $Y2=0.1350
r16 4 11 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2305 $Y2=0.1350
r17 4 19 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.2430 $Y=0.1350 $X2=0.2535 $Y2=0.1350
.ends

.subckt PM_AOI31xp67_ASAP7_75t_R%NET23 VSS 23 40 43 45 48 49 52 53 1 16 2 17 21
+ 3 18 4 19 5 20
c1 1 VSS 0.00807683f
c2 2 VSS 0.00681803f
c3 3 VSS 0.00543807f
c4 4 VSS 0.00970135f
c5 5 VSS 0.00989989f
c6 16 VSS 0.00369439f
c7 17 VSS 0.00335354f
c8 18 VSS 0.00228839f
c9 19 VSS 0.00459213f
c10 20 VSS 0.00450914f
c11 21 VSS 0.0439037f
r1 53 51 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r2 5 51 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5400 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r3 20 5 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.2025 $X2=0.5400 $Y2=0.2025
r4 52 20 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.2025 $X2=0.5255 $Y2=0.2025
r5 49 47 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r6 4 47 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r7 19 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r8 48 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r9 45 44 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r10 16 44 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r11 43 42 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r12 41 42 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1720 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r13 2 41 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1600 $Y=0.2025 $X2=0.1720 $Y2=0.2025
r14 17 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1600 $Y2=0.2025
r15 40 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r16 5 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.2025
+ $X2=0.5400 $Y2=0.2340
r17 4 35 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.2340
r18 1 31 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0520 $Y2=0.2340
r19 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r20 36 37 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.2340 $X2=0.5400 $Y2=0.2340
r21 35 36 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4860 $Y2=0.2340
r22 34 35 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.2340 $X2=0.4320 $Y2=0.2340
r23 33 34 18.8884 $w=1.3e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.3510 $Y2=0.2340
r24 32 33 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2315
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r25 28 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0610
+ $Y=0.2340 $X2=0.0790 $Y2=0.2340
r26 28 31 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0610
+ $Y=0.2340 $X2=0.0520 $Y2=0.2340
r27 27 29 5.13018 $w=1.3e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1010
+ $Y=0.2340 $X2=0.0790 $Y2=0.2340
r28 26 27 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1255
+ $Y=0.2340 $X2=0.1010 $Y2=0.2340
r29 25 32 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1865
+ $Y=0.2340 $X2=0.2315 $Y2=0.2340
r30 24 25 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1865 $Y2=0.2340
r31 21 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r32 21 26 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1255 $Y2=0.2340
r33 3 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.2340
r34 18 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2680 $Y2=0.2025
r35 23 18 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r36 1 16 1e-05
.ends

.subckt PM_AOI31xp67_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00408844f
.ends

.subckt PM_AOI31xp67_ASAP7_75t_R%NET29 VSS 12 13 28 29 1 7 9 2 8
c1 1 VSS 0.00971623f
c2 2 VSS 0.00468496f
c3 7 VSS 0.00452983f
c4 8 VSS 0.00229022f
c5 9 VSS 0.0325824f
r1 29 27 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r2 2 27 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0675 $X2=0.4320 $Y2=0.0675
r4 28 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4175 $Y2=0.0675
r5 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4320 $Y2=0.0360
r6 23 24 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3935
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r7 22 23 11.4263 $w=1.3e-08 $l=4.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.3445
+ $Y=0.0360 $X2=0.3935 $Y2=0.0360
r8 21 22 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3065
+ $Y=0.0360 $X2=0.3445 $Y2=0.0360
r9 20 21 8.51143 $w=1.3e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.3065 $Y2=0.0360
r10 19 20 10.0272 $w=1.3e-08 $l=4.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.2270
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r11 18 19 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1730
+ $Y=0.0360 $X2=0.2270 $Y2=0.0360
r12 17 18 9.91056 $w=1.3e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1305
+ $Y=0.0360 $X2=0.1730 $Y2=0.0360
r13 16 17 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1120
+ $Y=0.0360 $X2=0.1305 $Y2=0.0360
r14 14 16 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1030
+ $Y=0.0360 $X2=0.1120 $Y2=0.0360
r15 9 14 1.39914 $w=1.3e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.0970
+ $Y=0.0360 $X2=0.1030 $Y2=0.0360
r16 1 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1120 $Y2=0.0360
r17 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r18 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r19 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r20 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.0935 $Y2=0.0675
.ends

.subckt PM_AOI31xp67_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.0462333f
.ends

.subckt PM_AOI31xp67_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00657531f
.ends

.subckt PM_AOI31xp67_ASAP7_75t_R%NET30 VSS 15 29 30 32 1 2 11 13 10 3 12
c1 1 VSS 0.00368641f
c2 2 VSS 0.00337807f
c3 3 VSS 0.00304832f
c4 10 VSS 0.00296491f
c5 11 VSS 0.00222654f
c6 12 VSS 0.00240917f
c7 13 VSS 0.00285185f
r1 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.0675 $X2=0.5920 $Y2=0.0675
r2 32 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0675 $X2=0.5795 $Y2=0.0675
r3 30 28 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0675 $X2=0.5005 $Y2=0.0675
r4 2 28 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.0675 $X2=0.5005 $Y2=0.0675
r5 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0675 $X2=0.4860 $Y2=0.0675
r6 29 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4715 $Y2=0.0675
r7 3 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0675
+ $X2=0.5940 $Y2=0.0900
r8 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0675
+ $X2=0.4860 $Y2=0.0900
r9 24 25 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.5690
+ $Y=0.0900 $X2=0.5940 $Y2=0.0900
r10 23 24 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.5395
+ $Y=0.0900 $X2=0.5690 $Y2=0.0900
r11 22 23 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.5105
+ $Y=0.0900 $X2=0.5395 $Y2=0.0900
r12 21 22 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.0900 $X2=0.5105 $Y2=0.0900
r13 20 21 5.59655 $w=1.3e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.4620
+ $Y=0.0900 $X2=0.4860 $Y2=0.0900
r14 19 20 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4330
+ $Y=0.0900 $X2=0.4620 $Y2=0.0900
r15 18 19 6.99569 $w=1.3e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.4030
+ $Y=0.0900 $X2=0.4330 $Y2=0.0900
r16 17 18 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0900 $X2=0.4030 $Y2=0.0900
r17 13 17 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3665
+ $Y=0.0900 $X2=0.3780 $Y2=0.0900
r18 16 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.0945
+ $X2=0.3780 $Y2=0.0900
r19 1 16 23.8708 $w=2.02e-08 $l=4.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.3780 $Y=0.0540 $X2=0.3780 $Y2=0.0945
r20 15 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r21 10 14 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3800 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r22 1 10 1e-05
.ends

.subckt PM_AOI31xp67_ASAP7_75t_R%A1 VSS 20 3 4 1 5 6 7
c1 1 VSS 0.00403619f
c2 3 VSS 0.0427218f
c3 4 VSS 0.0424653f
c4 5 VSS 0.00735152f
c5 6 VSS 0.0121743f
c6 7 VSS 0.0116317f
c7 8 VSS 0.00449215f
r1 7 8 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6750 $Y=0.1665 $X2=0.6750 $Y2=0.1350
r2 6 8 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1125 $X2=0.6750 $Y2=0.1350
r3 8 24 1.26818 $w=1.72857e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6750 $Y=0.1350 $X2=0.6645 $Y2=0.1350
r4 23 24 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6355
+ $Y=0.1350 $X2=0.6645 $Y2=0.1350
r5 22 23 6.99569 $w=1.3e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.6055
+ $Y=0.1350 $X2=0.6355 $Y2=0.1350
r6 21 22 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.5895
+ $Y=0.1350 $X2=0.6055 $Y2=0.1350
r7 20 21 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5895 $Y2=0.1350
r8 20 5 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5555 $Y2=0.1350
r9 4 16 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1350
r10 20 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1350
+ $X2=0.5670 $Y2=0.1350
r11 15 16 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.5575
+ $Y=0.1350 $X2=0.5670 $Y2=0.1350
r12 13 15 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.5545 $Y=0.1350 $X2=0.5575 $Y2=0.1350
r13 12 13 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5400 $Y=0.1350 $X2=0.5545 $Y2=0.1350
r14 11 12 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5255 $Y=0.1350 $X2=0.5400 $Y2=0.1350
r15 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r16 1 10 3.20232 $w=2.13909e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5020 $Y2=0.1350
r17 1 11 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5255 $Y2=0.1350
r18 3 10 0.905388 $w=2.07755e-07 $l=1.1e-08 $layer=LIG $thickness=5.52727e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5020 $Y2=0.1350
r19 3 11 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5255 $Y2=0.1350
.ends

.subckt PM_AOI31xp67_ASAP7_75t_R%A2 VSS 19 3 4 1 7 6 5 8
c1 1 VSS 0.0109973f
c2 3 VSS 0.0466083f
c3 4 VSS 0.0461039f
c4 5 VSS 0.00430188f
c5 6 VSS 0.00528257f
c6 7 VSS 0.00439678f
c7 8 VSS 0.00468801f
r1 7 25 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0720 $X2=0.2970 $Y2=0.0900
r2 5 8 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1125 $X2=0.2970 $Y2=0.1350
r3 5 25 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1125 $X2=0.2970 $Y2=0.0900
r4 8 22 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1350 $X2=0.3155 $Y2=0.1350
r5 4 17 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1340
r6 21 22 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.3445
+ $Y=0.1350 $X2=0.3155 $Y2=0.1350
r7 19 6 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.3800 $Y2=0.1350
r8 6 21 8.27824 $w=1.3e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3800
+ $Y=0.1350 $X2=0.3445 $Y2=0.1350
r9 15 17 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4465 $Y=0.1340 $X2=0.4590 $Y2=0.1340
r10 14 15 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4320 $Y=0.1340 $X2=0.4465 $Y2=0.1340
r11 13 14 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4175 $Y=0.1340 $X2=0.4320 $Y2=0.1340
r12 11 13 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.4145 $Y=0.1340 $X2=0.4175 $Y2=0.1340
r13 10 11 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.4050
+ $Y=0.1340 $X2=0.4145 $Y2=0.1340
r14 19 10 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1340
r15 1 10 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.3955
+ $Y=0.1340 $X2=0.4050 $Y2=0.1340
r16 1 12 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.3955
+ $Y=0.1340 $X2=0.3945 $Y2=0.1340
r17 3 10 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4050 $Y2=0.1340
r18 3 12 0.610027 $w=2.16919e-07 $l=1.05475e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.4050 $Y=0.1350 $X2=0.3945 $Y2=0.1340
r19 3 13 1.79147 $w=1.8466e-07 $l=1.25399e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4175 $Y2=0.1340
.ends

.subckt PM_AOI31xp67_ASAP7_75t_R%Y VSS 31 26 47 50 67 68 2 21 22 1 13 16 15 17
+ 4 3 20 18 14 23 19 24
c1 1 VSS 0.00559539f
c2 2 VSS 0.00286645f
c3 3 VSS 0.00479122f
c4 4 VSS 0.0165118f
c5 13 VSS 0.00329753f
c6 14 VSS 0.0021398f
c7 15 VSS 0.00240953f
c8 16 VSS 0.000674098f
c9 17 VSS 0.00731234f
c10 18 VSS 0.0128917f
c11 19 VSS 0.000673989f
c12 20 VSS 0.00610522f
c13 21 VSS 0.000816538f
c14 22 VSS 0.000420816f
c15 23 VSS 0.000793832f
c16 24 VSS 0.00242386f
r1 68 66 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.0675 $X2=0.5545 $Y2=0.0675
r2 3 66 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5400 $Y=0.0675 $X2=0.5545 $Y2=0.0675
r3 14 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.0675 $X2=0.5400 $Y2=0.0675
r4 67 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.0675 $X2=0.5255 $Y2=0.0675
r5 3 63 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.0675
+ $X2=0.5400 $Y2=0.0360
r6 63 64 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.0360 $X2=0.5785 $Y2=0.0360
r7 18 60 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.6240
+ $Y=0.0360 $X2=0.6490 $Y2=0.0360
r8 18 64 10.6101 $w=1.3e-08 $l=4.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.6240
+ $Y=0.0360 $X2=0.5785 $Y2=0.0360
r9 58 59 23.8708 $w=2.02e-08 $l=4.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6490 $Y=0.0360 $X2=0.6490 $Y2=0.0765
r10 58 60 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6490 $Y=0.0360
+ $X2=0.6490 $Y2=0.0360
r11 57 59 22.9867 $w=2.02e-08 $l=3.9e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6490 $Y=0.1155 $X2=0.6490 $Y2=0.0765
r12 56 57 4.71523 $w=2.02e-08 $l=8e-09 $layer=LISD $thickness=2.7e-08 $X=0.6490
+ $Y=0.1235 $X2=0.6490 $Y2=0.1155
r13 55 56 6.77814 $w=2.02e-08 $l=1.15e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6490 $Y=0.1350 $X2=0.6490 $Y2=0.1235
r14 54 55 11.1987 $w=2.02e-08 $l=1.9e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6490 $Y=0.1540 $X2=0.6490 $Y2=0.1350
r15 4 53 23.8708 $w=2.02e-08 $l=4.05e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6490 $Y=0.1935 $X2=0.6490 $Y2=0.2340
r16 4 54 23.2814 $w=2.02e-08 $l=3.95e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.6490 $Y=0.1935 $X2=0.6490 $Y2=0.1540
r17 51 53 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6490 $Y=0.2340
+ $X2=0.6490 $Y2=0.2340
r18 20 51 6.41272 $w=1.3e-08 $l=2.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.6215
+ $Y=0.2340 $X2=0.6490 $Y2=0.2340
r19 20 24 4.76361 $w=1.46364e-08 $l=2.75e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6215 $Y=0.2340 $X2=0.5940 $Y2=0.2340
r20 19 45 2.45586 $w=1.44e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5940 $Y=0.2160 $X2=0.5940 $Y2=0.2035
r21 19 24 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.2160 $X2=0.5940 $Y2=0.2340
r22 50 49 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r23 48 49 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2260 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r24 2 48 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2140 $Y=0.2025 $X2=0.2260 $Y2=0.2025
r25 15 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2140 $Y2=0.2025
r26 47 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r27 23 45 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.1945 $X2=0.5940 $Y2=0.2035
r28 2 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.1980
r29 44 45 3.9716 $w=1.39211e-08 $l=2.51098e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5695 $Y=0.1980 $X2=0.5940 $Y2=0.2035
r30 43 44 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.5535
+ $Y=0.1980 $X2=0.5695 $Y2=0.1980
r31 42 43 15.7403 $w=1.3e-08 $l=6.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.1980 $X2=0.5535 $Y2=0.1980
r32 41 42 28.7989 $w=1.3e-08 $l=1.235e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.3625 $Y=0.1980 $X2=0.4860 $Y2=0.1980
r33 40 41 15.2739 $w=1.3e-08 $l=6.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1980 $X2=0.3625 $Y2=0.1980
r34 17 22 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2700 $Y=0.1980 $X2=0.2430 $Y2=0.1980
r35 17 40 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1980 $X2=0.2970 $Y2=0.1980
r36 37 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1980 $X2=0.2295 $Y2=0.1980
r37 22 35 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.1980 $X2=0.2430 $Y2=0.1765
r38 22 38 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.1980 $X2=0.2295 $Y2=0.1980
r39 34 35 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1540 $X2=0.2430 $Y2=0.1765
r40 33 34 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1540
r41 16 30 5.93557 $w=1.41538e-08 $l=3.15839e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.1035 $X2=0.2407 $Y2=0.0720
r42 16 33 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1035 $X2=0.2430 $Y2=0.1350
r43 31 30 0.739822 $w=1.8e-08 $l=7.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.2480
+ $Y=0.0720 $X2=0.2407 $Y2=0.0720
r44 29 30 1.73815 $w=1.6e-08 $l=1.12e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.0720 $X2=0.2407 $Y2=0.0720
r45 28 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0720 $X2=0.2295 $Y2=0.0720
r46 27 28 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2050
+ $Y=0.0720 $X2=0.2160 $Y2=0.0720
r47 21 27 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2025
+ $Y=0.0720 $X2=0.2050 $Y2=0.0720
r48 1 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0540
+ $X2=0.2160 $Y2=0.0720
r49 13 1 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0540 $X2=0.2140 $Y2=0.0540
r50 26 13 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0540 $X2=0.2015 $Y2=0.0540
.ends


*
.SUBCKT AOI31xp67_ASAP7_75t_R VSS VDD A3 B A2 A1 Y
*
* VSS VSS
* VDD VDD
* A3 A3
* B B
* A2 A2
* A1 A1
* Y Y
*
*

MM4 N_MM4_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@2 N_MM4@2_d N_MM4@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM7_g N_MM3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3@2 N_MM3@2_d N_MM7@2_g N_MM3@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM6_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2@2 N_MM2@2_d N_MM6@2_g N_MM2@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10@2 N_MM10@2_d N_MM4@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM5_g N_MM9_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9@2 N_MM9@2_d N_MM9@2_g N_MM9@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7@2 N_MM7@2_d N_MM7@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM6_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6@2 N_MM6@2_d N_MM6@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AOI31xp67_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AOI31xp67_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AOI31xp67_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_AOI31xp67_ASAP7_75t_R%noxref_12
cc_1 N_noxref_12_1 N_MM4_g 0.00221001f
cc_2 N_noxref_12_1 N_NET23_16 0.0360714f
cc_3 N_noxref_12_1 N_noxref_11_1 0.00177274f
x_PM_AOI31xp67_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_AOI31xp67_ASAP7_75t_R%noxref_14
cc_4 N_noxref_14_1 N_MM9@2_g 0.00152713f
cc_5 N_noxref_14_1 N_NET23_18 0.0358988f
cc_6 N_noxref_14_1 N_noxref_13_1 0.00138916f
x_PM_AOI31xp67_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_AOI31xp67_ASAP7_75t_R%noxref_16
cc_7 N_noxref_16_1 N_MM7_g 0.00159954f
cc_8 N_noxref_16_1 N_NET23_19 0.000668154f
cc_9 N_noxref_16_1 N_noxref_13_1 0.000477777f
cc_10 N_noxref_16_1 N_noxref_14_1 0.007665f
cc_11 N_noxref_16_1 N_noxref_15_1 0.00123f
x_PM_AOI31xp67_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_AOI31xp67_ASAP7_75t_R%noxref_11
cc_12 N_noxref_11_1 N_MM4_g 0.00228763f
cc_13 N_noxref_11_1 N_NET23_16 0.000477252f
x_PM_AOI31xp67_ASAP7_75t_R%A3 VSS A3 N_MM4_g N_MM4@2_g N_A3_7 N_A3_1 N_A3_10
+ PM_AOI31xp67_ASAP7_75t_R%A3
x_PM_AOI31xp67_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_AOI31xp67_ASAP7_75t_R%noxref_19
cc_14 N_noxref_19_1 N_MM6@2_g 0.000658581f
cc_15 N_noxref_19_1 N_Y_4 0.00456345f
cc_16 N_noxref_19_1 N_noxref_17_1 0.0080385f
cc_17 N_noxref_19_1 N_noxref_18_1 0.00198854f
x_PM_AOI31xp67_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_AOI31xp67_ASAP7_75t_R%noxref_18
cc_18 N_noxref_18_1 N_MM6@2_g 0.000665844f
cc_19 N_noxref_18_1 N_Y_4 0.00458151f
cc_20 N_noxref_18_1 N_noxref_17_1 0.00804671f
x_PM_AOI31xp67_ASAP7_75t_R%B VSS B N_MM5_g N_MM9@2_g N_B_8 N_B_5 N_B_6 N_B_10
+ N_B_1 N_B_9 N_B_7 PM_AOI31xp67_ASAP7_75t_R%B
cc_21 N_B_8 N_MM4@2_g 0.000560901f
cc_22 N_B_5 N_A3_7 0.000693988f
cc_23 N_B_6 N_A3_7 0.000720143f
cc_24 N_B_10 N_A3_1 0.00127368f
cc_25 N_B_10 N_A3_7 0.00186814f
cc_26 N_MM5_g N_MM4@2_g 0.0059152f
x_PM_AOI31xp67_ASAP7_75t_R%NET23 VSS N_MM9@2_s N_MM10@2_d N_MM9_s N_MM10_d
+ N_MM7_d N_MM7@2_d N_MM6_d N_MM6@2_d N_NET23_1 N_NET23_16 N_NET23_2 N_NET23_17
+ N_NET23_21 N_NET23_3 N_NET23_18 N_NET23_4 N_NET23_19 N_NET23_5 N_NET23_20
+ PM_AOI31xp67_ASAP7_75t_R%NET23
cc_27 N_NET23_1 N_MM4@2_g 0.00130793f
cc_28 N_NET23_16 N_MM4@2_g 0.000490744f
cc_29 N_NET23_2 N_MM4@2_g 0.000695186f
cc_30 N_NET23_17 N_A3_1 0.0015577f
cc_31 N_NET23_21 N_MM4@2_g 0.00164698f
cc_32 N_NET23_21 N_A3_10 0.00195422f
cc_33 N_NET23_1 N_MM4_g 0.00200906f
cc_34 N_NET23_16 N_MM4_g 0.0333552f
cc_35 N_NET23_17 N_MM4@2_g 0.0342072f
cc_36 N_NET23_2 N_MM9@2_g 0.000839165f
cc_37 N_NET23_17 N_MM9@2_g 0.000394869f
cc_38 N_NET23_3 N_MM9@2_g 0.000833663f
cc_39 N_NET23_2 N_MM5_g 0.00146825f
cc_40 N_NET23_18 N_B_1 0.00172273f
cc_41 N_NET23_21 N_MM9@2_g 0.00244601f
cc_42 N_NET23_21 N_B_9 0.00253235f
cc_43 N_NET23_17 N_MM5_g 0.0331307f
cc_44 N_NET23_18 N_MM9@2_g 0.0347356f
cc_45 N_NET23_4 N_MM7@2_g 0.00214826f
cc_46 N_NET23_3 N_MM7@2_g 0.000712458f
cc_47 N_NET23_19 N_A2_1 0.00193686f
cc_48 N_NET23_19 N_MM7_g 0.0183812f
cc_49 N_NET23_19 N_MM7@2_g 0.0497318f
cc_50 N_NET23_5 N_MM6@2_g 0.00185067f
cc_51 N_NET23_20 N_A1_1 0.00222344f
cc_52 N_NET23_20 N_MM6_g 0.0183527f
cc_53 N_NET23_20 N_MM6@2_g 0.0493815f
x_PM_AOI31xp67_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_AOI31xp67_ASAP7_75t_R%noxref_13
cc_54 N_noxref_13_1 N_MM9@2_g 0.00890749f
cc_55 N_noxref_13_1 N_MM7_g 0.00075126f
cc_56 N_noxref_13_1 N_NET23_18 0.000496275f
cc_57 N_noxref_13_1 N_NET29_9 0.000291841f
cc_58 N_noxref_13_1 N_NET30_10 0.000646426f
cc_59 N_noxref_13_1 N_Y_13 0.000743044f
x_PM_AOI31xp67_ASAP7_75t_R%NET29 VSS N_MM4_d N_MM4@2_d N_MM3_s N_MM3@2_s
+ N_NET29_1 N_NET29_7 N_NET29_9 N_NET29_2 N_NET29_8
+ PM_AOI31xp67_ASAP7_75t_R%NET29
cc_60 N_NET29_1 N_MM4@2_g 0.00197873f
cc_61 N_NET29_7 N_A3_1 0.00204582f
cc_62 N_NET29_7 N_MM4_g 0.0182808f
cc_63 N_NET29_7 N_MM4@2_g 0.050442f
cc_64 N_NET29_9 N_B_8 0.00234078f
cc_65 N_NET29_9 N_MM9@2_g 0.00435002f
cc_66 N_NET29_2 N_MM7@2_g 0.00178562f
cc_67 N_NET29_8 N_A2_1 0.0020807f
cc_68 N_NET29_9 N_A2_7 0.00475644f
cc_69 N_NET29_8 N_MM7_g 0.0182772f
cc_70 N_NET29_8 N_MM7@2_g 0.0495034f
x_PM_AOI31xp67_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_AOI31xp67_ASAP7_75t_R%noxref_17
cc_71 N_noxref_17_1 N_MM6@2_g 0.00371316f
cc_72 N_noxref_17_1 N_NET30_12 0.0363043f
cc_73 N_noxref_17_1 N_Y_4 0.00690334f
x_PM_AOI31xp67_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_AOI31xp67_ASAP7_75t_R%noxref_15
cc_74 N_noxref_15_1 N_MM7_g 0.0017298f
cc_75 N_noxref_15_1 N_NET30_10 0.0360377f
cc_76 N_noxref_15_1 N_noxref_13_1 0.0078498f
x_PM_AOI31xp67_ASAP7_75t_R%NET30 VSS N_MM3_d N_MM3@2_d N_MM2_s N_MM2@2_s
+ N_NET30_1 N_NET30_2 N_NET30_11 N_NET30_13 N_NET30_10 N_NET30_3 N_NET30_12
+ PM_AOI31xp67_ASAP7_75t_R%NET30
cc_77 N_NET30_1 N_A2_1 0.000596371f
cc_78 N_NET30_1 N_A2_6 0.000612158f
cc_79 N_NET30_2 N_MM7@2_g 0.00070839f
cc_80 N_NET30_1 N_MM7_g 0.00124065f
cc_81 N_NET30_11 N_A2_1 0.0019732f
cc_82 N_NET30_13 N_A2_6 0.00249384f
cc_83 N_NET30_13 N_A2_1 0.00294659f
cc_84 N_NET30_11 N_MM7@2_g 0.0331881f
cc_85 N_NET30_10 N_MM7_g 0.0353007f
cc_86 N_NET30_3 N_MM6@2_g 0.00154597f
cc_87 N_NET30_2 N_MM6_g 0.000732495f
cc_88 N_NET30_12 N_A1_1 0.00218081f
cc_89 N_NET30_13 N_A1_5 0.00229435f
cc_90 N_NET30_13 N_A1_1 0.00281931f
cc_91 N_NET30_11 N_MM6_g 0.0332828f
cc_92 N_NET30_12 N_MM6@2_g 0.0353598f
cc_93 N_NET30_13 N_NET29_8 0.00059447f
cc_94 N_NET30_2 N_NET29_2 0.00508278f
cc_95 N_NET30_11 N_NET29_8 0.00112154f
cc_96 N_NET30_1 N_NET29_2 0.00189294f
cc_97 N_NET30_13 N_NET29_9 0.00726951f
x_PM_AOI31xp67_ASAP7_75t_R%A1 VSS A1 N_MM6_g N_MM6@2_g N_A1_1 N_A1_5 N_A1_6
+ N_A1_7 PM_AOI31xp67_ASAP7_75t_R%A1
cc_98 N_MM6_g N_MM7@2_g 0.00457224f
x_PM_AOI31xp67_ASAP7_75t_R%A2 VSS A2 N_MM7_g N_MM7@2_g N_A2_1 N_A2_7 N_A2_6
+ N_A2_5 N_A2_8 PM_AOI31xp67_ASAP7_75t_R%A2
x_PM_AOI31xp67_ASAP7_75t_R%Y VSS Y N_MM5_d N_MM9_d N_MM9@2_d N_MM2_d N_MM2@2_d
+ N_Y_2 N_Y_21 N_Y_22 N_Y_1 N_Y_13 N_Y_16 N_Y_15 N_Y_17 N_Y_4 N_Y_3 N_Y_20
+ N_Y_18 N_Y_14 N_Y_23 N_Y_19 N_Y_24 PM_AOI31xp67_ASAP7_75t_R%Y
cc_99 N_Y_2 N_MM9@2_g 0.00204303f
cc_100 N_Y_21 N_MM9@2_g 0.000809466f
cc_101 N_Y_22 N_MM9@2_g 0.000757348f
cc_102 N_Y_1 N_MM9@2_g 0.00142535f
cc_103 N_Y_2 N_B_1 0.000645528f
cc_104 N_Y_13 N_MM5_g 0.00871502f
cc_105 N_Y_16 N_B_7 0.00343262f
cc_106 N_Y_15 N_B_1 0.00389109f
cc_107 N_Y_13 N_MM9@2_g 0.014688f
cc_108 N_Y_15 N_MM5_g 0.0318156f
cc_109 N_Y_15 N_MM9@2_g 0.0635972f
cc_110 N_Y_21 N_A2_6 0.000805472f
cc_111 N_Y_16 N_A2_5 0.00103451f
cc_112 N_Y_17 N_A2_8 0.00155218f
cc_113 N_Y_16 N_A2_8 0.0022071f
cc_114 N_Y_17 N_A2_6 0.00579974f
cc_115 N_Y_4 N_MM6@2_g 0.000629579f
cc_116 N_Y_3 N_MM6@2_g 0.00222381f
cc_117 N_Y_20 N_MM6@2_g 0.000797934f
cc_118 N_Y_18 N_A1_6 0.000979912f
cc_119 N_Y_17 N_A1_1 0.00113807f
cc_120 N_Y_4 N_A1_6 0.00174736f
cc_121 N_Y_4 N_A1_7 0.00182813f
cc_122 N_Y_14 N_A1_1 0.00268467f
cc_123 N_Y_4 N_A1_5 0.00287227f
cc_124 N_Y_23 N_A1_5 0.00302876f
cc_125 N_Y_14 N_MM6_g 0.018483f
cc_126 N_Y_14 N_MM6@2_g 0.0496668f
cc_127 N_Y_19 N_NET23_21 0.000161059f
cc_128 N_Y_2 N_NET23_21 0.000909366f
cc_129 N_Y_24 N_NET23_21 0.000329532f
cc_130 N_Y_17 N_NET23_4 0.00122194f
cc_131 N_Y_16 N_NET23_3 0.000508614f
cc_132 N_Y_15 N_NET23_17 0.000562552f
cc_133 N_Y_17 N_NET23_5 0.00142222f
cc_134 N_Y_17 N_NET23_3 0.000613924f
cc_135 N_Y_15 N_NET23_18 0.00174961f
cc_136 N_Y_2 N_NET23_2 0.00138315f
cc_137 N_Y_22 N_NET23_21 0.00218735f
cc_138 N_Y_2 N_NET23_3 0.00510943f
cc_139 N_Y_17 N_NET23_21 0.0267283f
cc_140 N_Y_16 N_NET29_9 0.000260458f
cc_141 N_Y_1 N_NET29_9 0.000914742f
cc_142 N_Y_21 N_NET29_9 0.00660877f
cc_143 N_Y_4 N_NET30_13 0.000206169f
cc_144 N_Y_3 N_NET30_13 0.000856257f
cc_145 N_Y_14 N_NET30_13 0.000566575f
cc_146 N_Y_3 N_NET30_3 0.00689012f
cc_147 N_Y_17 N_NET30_13 0.000738005f
cc_148 N_Y_14 N_NET30_12 0.00218825f
cc_149 N_Y_3 N_NET30_2 0.00135936f
cc_150 N_Y_4 N_NET30_12 0.00205357f
cc_151 N_Y_18 N_NET30_13 0.00701629f
*END of AOI31xp67_ASAP7_75t_R.pxi
.ENDS
** Design:	AOI321xp33_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AOI321xp33_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AOI321xp33_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AOI321xp33_ASAP7_75t_R%NET026 VSS 2 3 1
c1 1 VSS 0.00085891f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0540 $X2=0.3240 $Y2=0.0540
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0540 $X2=0.3240 $Y2=0.0540
.ends

.subckt PM_AOI321xp33_ASAP7_75t_R%NET30 VSS 2 3 1
c1 1 VSS 0.000941975f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_AOI321xp33_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.0424523f
.ends

.subckt PM_AOI321xp33_ASAP7_75t_R%NET29 VSS 2 3 1
c1 1 VSS 0.00094051f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_AOI321xp33_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.0425023f
.ends

.subckt PM_AOI321xp33_ASAP7_75t_R%NET23 VSS 12 13 24 27 7 1 9 2 8
c1 1 VSS 0.00862637f
c2 2 VSS 0.00615459f
c3 7 VSS 0.00449525f
c4 8 VSS 0.00342683f
c5 9 VSS 0.00687895f
r1 27 26 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r2 25 26 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2260 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r3 2 25 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2140 $Y=0.2025 $X2=0.2260 $Y2=0.2025
r4 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2140 $Y2=0.2025
r5 24 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r6 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.1980
r7 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2025
+ $Y=0.1980 $X2=0.2160 $Y2=0.1980
r8 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1980 $X2=0.2025 $Y2=0.1980
r9 18 19 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.1980 $X2=0.1890 $Y2=0.1980
r10 17 18 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1980 $X2=0.1620 $Y2=0.1980
r11 16 17 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1215
+ $Y=0.1980 $X2=0.1350 $Y2=0.1980
r12 15 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.1980 $X2=0.1215 $Y2=0.1980
r13 14 15 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0970
+ $Y=0.1980 $X2=0.1080 $Y2=0.1980
r14 9 14 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.1980 $X2=0.0970 $Y2=0.1980
r15 1 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.1980
r16 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r17 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r18 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r19 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
.ends

.subckt PM_AOI321xp33_ASAP7_75t_R%A3 VSS 9 3 1 6
c1 1 VSS 0.00481294f
c2 3 VSS 0.0820804f
c3 4 VSS 0.011835f
c4 5 VSS 0.0116426f
c5 6 VSS 0.00313729f
c6 7 VSS 0.00187052f
r1 5 7 3.2503 $w=1.53684e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1540 $X2=0.0270 $Y2=0.1350
r2 4 7 11.6451 $w=1.38182e-08 $l=5.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0800 $X2=0.0270 $Y2=0.1350
r3 9 6 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0540 $Y2=0.1350
r4 6 7 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.1350 $X2=0.0270 $Y2=0.1350
r5 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r6 9 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AOI321xp33_ASAP7_75t_R%B1 VSS 6 3 1 4
c1 1 VSS 0.00557387f
c2 3 VSS 0.0353407f
c3 4 VSS 0.00424541f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.0980
r2 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_AOI321xp33_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.00554638f
.ends

.subckt PM_AOI321xp33_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.00473487f
.ends

.subckt PM_AOI321xp33_ASAP7_75t_R%A2 VSS 4 3 1
c1 1 VSS 0.00684384f
c2 3 VSS 0.0466603f
c3 4 VSS 0.00800407f
r1 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r2 4 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AOI321xp33_ASAP7_75t_R%C VSS 6 3 4 1
c1 1 VSS 0.0074095f
c2 3 VSS 0.035258f
c3 4 VSS 0.00515471f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.0980
r2 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AOI321xp33_ASAP7_75t_R%A1 VSS 6 3 1 4
c1 1 VSS 0.00833305f
c2 3 VSS 0.0462427f
c3 4 VSS 0.00485879f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.0980
r2 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AOI321xp33_ASAP7_75t_R%B2 VSS 6 3 1 4
c1 1 VSS 0.00640274f
c2 3 VSS 0.00835705f
c3 4 VSS 0.00408339f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.0980
r2 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
.ends

.subckt PM_AOI321xp33_ASAP7_75t_R%Y VSS 33 22 23 47 54 55 15 10 1 11 16 14 2 3
+ 12 17 19
c1 1 VSS 0.00785409f
c2 2 VSS 0.00297509f
c3 3 VSS 0.00545643f
c4 10 VSS 0.00313767f
c5 11 VSS 0.000398848f
c6 12 VSS 0.00255416f
c7 13 VSS 6.0498e-20
c8 14 VSS 0.00213954f
c9 15 VSS 0.0187545f
c10 16 VSS 0.000769627f
c11 17 VSS 0.00210799f
c12 18 VSS 0.00277642f
c13 19 VSS 0.000735372f
r1 55 53 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r2 2 53 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r3 14 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r4 54 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r5 2 50 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.1980
r6 50 51 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1980 $X2=0.3375 $Y2=0.1980
r7 48 51 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1980 $X2=0.3375 $Y2=0.1980
r8 16 19 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3780 $Y=0.1980 $X2=0.4050 $Y2=0.1980
r9 16 48 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.1980 $X2=0.3510 $Y2=0.1980
r10 19 45 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.1980 $X2=0.4050 $Y2=0.1765
r11 12 3 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.0540 $X2=0.3760 $Y2=0.0540
r12 47 12 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0540 $X2=0.3635 $Y2=0.0540
r13 44 45 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1170 $X2=0.4050 $Y2=0.1765
r14 17 18 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.0575 $X2=0.4050 $Y2=0.0360
r15 17 44 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0575 $X2=0.4050 $Y2=0.1170
r16 3 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.0540
+ $X2=0.3780 $Y2=0.0360
r17 18 43 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.0360 $X2=0.3915 $Y2=0.0360
r18 42 43 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0360 $X2=0.3915 $Y2=0.0360
r19 41 42 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3645
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r20 40 41 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0360 $X2=0.3645 $Y2=0.0360
r21 39 40 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3260
+ $Y=0.0360 $X2=0.3510 $Y2=0.0360
r22 38 39 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3080
+ $Y=0.0360 $X2=0.3260 $Y2=0.0360
r23 37 38 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.3080 $Y2=0.0360
r24 36 37 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2720
+ $Y=0.0360 $X2=0.2970 $Y2=0.0360
r25 35 36 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2540
+ $Y=0.0360 $X2=0.2720 $Y2=0.0360
r26 34 35 0.874462 $w=1.3e-08 $l=3.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.2502
+ $Y=0.0360 $X2=0.2540 $Y2=0.0360
r27 33 34 0.524677 $w=1.3e-08 $l=2.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.2480
+ $Y=0.0360 $X2=0.2502 $Y2=0.0360
r28 33 32 1.69063 $w=1.3e-08 $l=7.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.2480
+ $Y=0.0360 $X2=0.2407 $Y2=0.0360
r29 31 32 2.04041 $w=1.3e-08 $l=8.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.2320
+ $Y=0.0360 $X2=0.2407 $Y2=0.0360
r30 30 31 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2275
+ $Y=0.0360 $X2=0.2320 $Y2=0.0360
r31 29 30 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.2275 $Y2=0.0360
r32 15 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2025
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r33 11 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0945 $X2=0.2140 $Y2=0.0945
r34 1 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0540
+ $X2=0.2160 $Y2=0.0360
r35 25 26 0.264706 $w=1.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2260 $Y=0.0725 $X2=0.2305 $Y2=0.0725
r36 1 25 0.705882 $w=1.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2140 $Y=0.0725 $X2=0.2260 $Y2=0.0725
r37 13 1 0.735294 $w=1.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0725 $X2=0.2140 $Y2=0.0725
r38 23 21 0.0675676 $w=3.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0455 $X2=0.2305 $Y2=0.0455
r39 1 21 0.391892 $w=3.7e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.0455 $X2=0.2305 $Y2=0.0455
r40 1 26 0.471383 $w=3.35517e-08 $l=3.06472e-08 $layer=N_src_drn
+ $thickness=1e-09 $X=0.2160 $Y=0.0455 $X2=0.2305 $Y2=0.0725
r41 10 1 0.391892 $w=3.7e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0455 $X2=0.2160 $Y2=0.0455
r42 22 10 0.0675676 $w=3.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0455 $X2=0.2015 $Y2=0.0455
.ends

.subckt PM_AOI321xp33_ASAP7_75t_R%NET013 VSS 12 13 22 7 1 8 2 9
c1 1 VSS 0.00492126f
c2 2 VSS 0.00511764f
c3 7 VSS 0.00218907f
c4 8 VSS 0.00225542f
c5 9 VSS 0.0131763f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3760 $Y2=0.2025
r2 22 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r3 2 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.2340
r4 18 19 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3395
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r5 17 18 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3080
+ $Y=0.2340 $X2=0.3395 $Y2=0.2340
r6 16 17 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.2340 $X2=0.3080 $Y2=0.2340
r7 15 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2835
+ $Y=0.2340 $X2=0.2970 $Y2=0.2340
r8 14 15 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.2835 $Y2=0.2340
r9 9 14 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2585
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r10 1 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.2340
r11 12 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r12 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r13 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r14 13 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
.ends


*
.SUBCKT AOI321xp33_ASAP7_75t_R VSS VDD A3 A2 A1 C B1 B2 Y
*
* VSS VSS
* VDD VDD
* A3 A3
* A2 A2
* A1 A1
* C C
* B1 B1
* B2 B2
* Y Y
*
*

MM4 N_MM4_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g N_MM3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM0_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM9_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM11 N_MM11_d N_MM8_g N_MM11_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM10 N_MM10_d N_MM4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM12 N_MM12_d N_MM0_g N_MM12_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM8_g N_MM8_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AOI321xp33_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AOI321xp33_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AOI321xp33_ASAP7_75t_R%NET026 VSS N_MM5_d N_MM11_s N_NET026_1
+ PM_AOI321xp33_ASAP7_75t_R%NET026
cc_1 N_NET026_1 N_MM9_g 0.0126998f
cc_2 N_NET026_1 N_MM8_g 0.0126111f
x_PM_AOI321xp33_ASAP7_75t_R%NET30 VSS N_MM3_d N_MM2_s N_NET30_1
+ PM_AOI321xp33_ASAP7_75t_R%NET30
cc_3 N_NET30_1 N_MM3_g 0.0172839f
cc_4 N_NET30_1 N_MM2_g 0.0171487f
x_PM_AOI321xp33_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_AOI321xp33_ASAP7_75t_R%noxref_15
cc_5 N_noxref_15_1 N_MM4_g 0.00221934f
x_PM_AOI321xp33_ASAP7_75t_R%NET29 VSS N_MM4_d N_MM3_s N_NET29_1
+ PM_AOI321xp33_ASAP7_75t_R%NET29
cc_6 N_NET29_1 N_MM4_g 0.0173543f
cc_7 N_NET29_1 N_MM3_g 0.0172743f
x_PM_AOI321xp33_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_AOI321xp33_ASAP7_75t_R%noxref_16
cc_8 N_noxref_16_1 N_MM4_g 0.00221256f
cc_9 N_noxref_16_1 N_noxref_15_1 0.00176928f
x_PM_AOI321xp33_ASAP7_75t_R%NET23 VSS N_MM10_d N_MM7_d N_MM6_d N_MM12_s
+ N_NET23_7 N_NET23_1 N_NET23_9 N_NET23_2 N_NET23_8
+ PM_AOI321xp33_ASAP7_75t_R%NET23
cc_10 N_NET23_7 N_A3_1 0.000685029f
cc_11 N_NET23_1 N_MM4_g 0.000939786f
cc_12 N_NET23_9 N_A3_6 0.00128131f
cc_13 N_NET23_7 N_MM4_g 0.034145f
cc_14 N_NET23_7 N_A2_1 0.00079996f
cc_15 N_NET23_1 N_MM3_g 0.000879863f
cc_16 N_NET23_9 N_A2 0.00118443f
cc_17 N_NET23_1 N_A2 0.0012945f
cc_18 N_NET23_7 N_MM3_g 0.0335084f
cc_19 N_NET23_2 N_MM2_g 0.000873416f
cc_20 N_NET23_9 N_A1_4 0.00112697f
cc_21 N_NET23_2 N_A1_4 0.00129672f
cc_22 N_NET23_8 N_MM2_g 0.0342621f
cc_23 N_NET23_8 N_C_1 0.000744697f
cc_24 N_NET23_2 N_C_4 0.000840829f
cc_25 N_NET23_2 N_MM0_g 0.000888931f
cc_26 N_NET23_8 N_MM0_g 0.0337964f
x_PM_AOI321xp33_ASAP7_75t_R%A3 VSS A3 N_MM4_g N_A3_1 N_A3_6
+ PM_AOI321xp33_ASAP7_75t_R%A3
x_PM_AOI321xp33_ASAP7_75t_R%B1 VSS B1 N_MM9_g N_B1_1 N_B1_4
+ PM_AOI321xp33_ASAP7_75t_R%B1
cc_27 N_B1_1 N_C_1 0.00116455f
cc_28 N_B1_4 N_C_4 0.00367739f
cc_29 N_MM9_g N_MM0_g 0.00625031f
x_PM_AOI321xp33_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_AOI321xp33_ASAP7_75t_R%noxref_18
cc_30 N_noxref_18_1 N_MM8_g 0.00159541f
cc_31 N_noxref_18_1 N_NET013_8 0.0364877f
cc_32 N_noxref_18_1 N_Y_14 0.000863584f
cc_33 N_noxref_18_1 N_noxref_17_1 0.00189902f
x_PM_AOI321xp33_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_AOI321xp33_ASAP7_75t_R%noxref_17
cc_34 N_noxref_17_1 N_MM8_g 0.00349598f
cc_35 N_noxref_17_1 N_NET013_8 0.000590033f
cc_36 N_noxref_17_1 N_Y_12 0.0278837f
x_PM_AOI321xp33_ASAP7_75t_R%A2 VSS A2 N_MM3_g N_A2_1
+ PM_AOI321xp33_ASAP7_75t_R%A2
cc_37 N_A2_1 N_MM4_g 0.0006597f
cc_38 N_A2_1 N_A3_1 0.00130265f
cc_39 N_A2 N_A3_6 0.00265118f
cc_40 N_MM3_g N_MM4_g 0.00611045f
x_PM_AOI321xp33_ASAP7_75t_R%C VSS C N_MM0_g N_C_4 N_C_1
+ PM_AOI321xp33_ASAP7_75t_R%C
cc_41 N_MM0_g N_MM2_g 0.00329319f
cc_42 N_C_4 N_A1_4 0.0049527f
x_PM_AOI321xp33_ASAP7_75t_R%A1 VSS A1 N_MM2_g N_A1_1 N_A1_4
+ PM_AOI321xp33_ASAP7_75t_R%A1
cc_43 N_A1_1 N_A2_1 0.00121341f
cc_44 N_A1_4 N_A2 0.00393573f
cc_45 N_MM2_g N_MM3_g 0.00615078f
x_PM_AOI321xp33_ASAP7_75t_R%B2 VSS B2 N_MM8_g N_B2_1 N_B2_4
+ PM_AOI321xp33_ASAP7_75t_R%B2
cc_46 N_B2_1 N_B1_1 0.00130341f
cc_47 N_B2_4 N_B1_4 0.00340374f
cc_48 N_MM8_g N_MM9_g 0.00757165f
x_PM_AOI321xp33_ASAP7_75t_R%Y VSS Y N_MM2_d N_MM0_d N_MM11_d N_MM9_d N_MM8_d
+ N_Y_15 N_Y_10 N_Y_1 N_Y_11 N_Y_16 N_Y_14 N_Y_2 N_Y_3 N_Y_12 N_Y_17 N_Y_19
+ PM_AOI321xp33_ASAP7_75t_R%Y
cc_49 N_Y_15 N_A2 0.00161937f
cc_50 N_Y_15 N_MM2_g 0.000641302f
cc_51 N_Y_10 N_A1_1 0.000647573f
cc_52 N_Y_1 N_A1_4 0.00132276f
cc_53 N_Y_1 N_MM2_g 0.00152282f
cc_54 N_Y_10 N_MM2_g 0.00981004f
cc_55 N_Y_11 N_MM2_g 0.0248709f
cc_56 N_Y_15 N_C_4 0.00113494f
cc_57 N_Y_1 N_MM0_g 0.00127804f
cc_58 N_Y_1 N_C_4 0.0018474f
cc_59 N_Y_11 N_MM0_g 0.005217f
cc_60 N_Y_10 N_MM0_g 0.0306992f
cc_61 N_Y_16 N_B1_4 0.000570438f
cc_62 N_Y_14 N_B1_1 0.000815217f
cc_63 N_Y_2 N_MM9_g 0.000919549f
cc_64 N_Y_15 N_B1_4 0.00137688f
cc_65 N_Y_2 N_B1_4 0.00215366f
cc_66 N_Y_14 N_MM9_g 0.0356016f
cc_67 N_Y_2 N_B2_1 0.000697718f
cc_68 N_Y_2 N_MM8_g 0.000899074f
cc_69 N_Y_3 N_MM8_g 0.000933765f
cc_70 N_Y_16 N_B2_4 0.00109994f
cc_71 N_Y_14 N_B2_1 0.00119684f
cc_72 N_Y_15 N_B2_4 0.00120568f
cc_73 N_Y_12 N_MM8_g 0.0109422f
cc_74 N_Y_17 N_B2_4 0.00654921f
cc_75 N_Y_14 N_MM8_g 0.0487869f
cc_76 N_Y_16 N_NET013_2 0.000633418f
cc_77 N_Y_19 N_NET013_9 0.000676724f
cc_78 N_Y_14 N_NET013_8 0.000714362f
cc_79 N_Y_17 N_NET013_2 0.000720076f
cc_80 N_Y_2 N_NET013_9 0.00096803f
cc_81 N_Y_14 N_NET013_7 0.00112742f
cc_82 N_Y_2 N_NET013_2 0.00242734f
cc_83 N_Y_2 N_NET013_1 0.00418801f
cc_84 N_Y_16 N_NET013_9 0.00931193f
x_PM_AOI321xp33_ASAP7_75t_R%NET013 VSS N_MM9_s N_MM12_d N_MM8_s N_NET013_7
+ N_NET013_1 N_NET013_8 N_NET013_2 N_NET013_9 PM_AOI321xp33_ASAP7_75t_R%NET013
cc_85 N_NET013_7 N_C_1 0.000734666f
cc_86 N_NET013_1 N_MM0_g 0.00094989f
cc_87 N_NET013_7 N_MM0_g 0.0346173f
cc_88 N_NET013_7 N_B1_1 0.000664781f
cc_89 N_NET013_1 N_MM9_g 0.00095181f
cc_90 N_NET013_7 N_MM9_g 0.0347767f
cc_91 N_NET013_8 N_B2_1 0.0007277f
cc_92 N_NET013_2 N_MM8_g 0.00106064f
cc_93 N_NET013_8 N_MM8_g 0.03486f
cc_94 N_NET013_7 N_NET23_2 0.00055449f
cc_95 N_NET013_9 N_NET23_9 0.00109119f
cc_96 N_NET013_1 N_NET23_2 0.00389832f
*END of AOI321xp33_ASAP7_75t_R.pxi
.ENDS
** Design:	AOI322xp5_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AOI322xp5_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AOI322xp5_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AOI322xp5_ASAP7_75t_R%NET52 VSS 2 3 1
c1 1 VSS 0.000962086f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2700 $Y2=0.0675
.ends

.subckt PM_AOI322xp5_ASAP7_75t_R%NET51 VSS 2 3 1
c1 1 VSS 0.000879498f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0540 $X2=0.1080 $Y2=0.0540
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0540 $X2=0.1080 $Y2=0.0540
.ends

.subckt PM_AOI322xp5_ASAP7_75t_R%NET50 VSS 2 3 1
c1 1 VSS 0.000875344f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0540 $X2=0.3780 $Y2=0.0540
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0540 $X2=0.3780 $Y2=0.0540
.ends

.subckt PM_AOI322xp5_ASAP7_75t_R%NET49 VSS 2 3 1
c1 1 VSS 0.000970332f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2160 $Y2=0.0675
.ends

.subckt PM_AOI322xp5_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.00624108f
.ends

.subckt PM_AOI322xp5_ASAP7_75t_R%B2 VSS 6 3 1 4
c1 1 VSS 0.00347696f
c2 3 VSS 0.0715143f
c3 4 VSS 0.014569f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.0980
r2 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AOI322xp5_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.0320247f
.ends

.subckt PM_AOI322xp5_ASAP7_75t_R%B1 VSS 6 3 1 4
c1 1 VSS 0.00699742f
c2 3 VSS 0.0458546f
c3 4 VSS 0.00413785f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.0980
r2 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AOI322xp5_ASAP7_75t_R%A3 VSS 6 3 1 4
c1 1 VSS 0.00771582f
c2 3 VSS 0.0466068f
c3 4 VSS 0.00492911f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.0980
r2 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_AOI322xp5_ASAP7_75t_R%C2 VSS 6 3 4 1
c1 1 VSS 0.00677128f
c2 3 VSS 0.0462891f
c3 4 VSS 0.00463114f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.0980
r2 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
.ends

.subckt PM_AOI322xp5_ASAP7_75t_R%A2 VSS 6 3 1 4
c1 1 VSS 0.00688477f
c2 3 VSS 0.00958784f
c3 4 VSS 0.00456113f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.0980
r2 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AOI322xp5_ASAP7_75t_R%A1 VSS 6 3 1 4
c1 1 VSS 0.0077695f
c2 3 VSS 0.00908874f
c3 4 VSS 0.00493039f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.0980
r2 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AOI322xp5_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.00473642f
.ends

.subckt PM_AOI322xp5_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.00573112f
.ends

.subckt PM_AOI322xp5_ASAP7_75t_R%NET27 VSS 16 17 35 38 40 10 1 13 11 2 12 3
c1 1 VSS 0.00722521f
c2 2 VSS 0.00603818f
c3 3 VSS 0.00314675f
c4 10 VSS 0.00353547f
c5 11 VSS 0.00337942f
c6 12 VSS 0.00216827f
c7 13 VSS 0.00753552f
r1 40 39 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r2 10 39 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r3 38 37 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r4 2 37 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1640 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r5 34 2 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1520 $Y=0.2025 $X2=0.1640 $Y2=0.2025
r6 11 34 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1520 $Y2=0.2025
r7 35 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r8 1 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.1980
r9 2 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.1980
r10 32 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.1980 $X2=0.0675 $Y2=0.1980
r11 30 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1980 $X2=0.0675 $Y2=0.1980
r12 29 30 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.1980 $X2=0.0810 $Y2=0.1980
r13 28 29 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1980 $X2=0.1080 $Y2=0.1980
r14 27 28 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1455
+ $Y=0.1980 $X2=0.1350 $Y2=0.1980
r15 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.1980 $X2=0.1755 $Y2=0.1980
r16 24 25 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1500
+ $Y=0.1980 $X2=0.1620 $Y2=0.1980
r17 24 27 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1500
+ $Y=0.1980 $X2=0.1455 $Y2=0.1980
r18 23 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1980 $X2=0.1755 $Y2=0.1980
r19 22 23 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2000
+ $Y=0.1980 $X2=0.1890 $Y2=0.1980
r20 21 22 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2180
+ $Y=0.1980 $X2=0.2000 $Y2=0.1980
r21 20 21 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1980 $X2=0.2180 $Y2=0.1980
r22 13 18 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.1980 $X2=0.2700 $Y2=0.1980
r23 13 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.1980 $X2=0.2430 $Y2=0.1980
r24 3 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.1980
r25 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r26 3 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r27 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r28 16 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r29 1 10 1e-05
.ends

.subckt PM_AOI322xp5_ASAP7_75t_R%C1 VSS 6 3 1 4
c1 1 VSS 0.00680149f
c2 3 VSS 0.00857902f
c3 4 VSS 0.004326f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.0980
r2 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
.ends

.subckt PM_AOI322xp5_ASAP7_75t_R%Y VSS 34 22 23 51 58 59 15 10 1 11 16 14 2 3
+ 12 17 19
c1 1 VSS 0.00643939f
c2 2 VSS 0.00281012f
c3 3 VSS 0.00553461f
c4 10 VSS 0.00282618f
c5 11 VSS 0.000465698f
c6 12 VSS 0.00259261f
c7 13 VSS 7.04036e-20
c8 14 VSS 0.00214559f
c9 15 VSS 0.0284543f
c10 16 VSS 0.000711061f
c11 17 VSS 0.00206266f
c12 18 VSS 0.00277543f
c13 19 VSS 0.000741384f
r1 59 57 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r2 2 57 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r3 14 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3780 $Y2=0.2025
r4 58 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r5 2 54 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.1980
r6 54 55 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.1980 $X2=0.3915 $Y2=0.1980
r7 52 55 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1980 $X2=0.3915 $Y2=0.1980
r8 16 19 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4320 $Y=0.1980 $X2=0.4590 $Y2=0.1980
r9 16 52 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.1980 $X2=0.4050 $Y2=0.1980
r10 19 49 3.24787 $w=1.72e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1980 $X2=0.4590 $Y2=0.1770
r11 12 3 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0540 $X2=0.4300 $Y2=0.0540
r12 51 12 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0540 $X2=0.4175 $Y2=0.0540
r13 48 49 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1645 $X2=0.4590 $Y2=0.1770
r14 47 48 11.0765 $w=1.3e-08 $l=4.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1170 $X2=0.4590 $Y2=0.1645
r15 17 18 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0575 $X2=0.4590 $Y2=0.0360
r16 17 47 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0575 $X2=0.4590 $Y2=0.1170
r17 3 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0540
+ $X2=0.4320 $Y2=0.0360
r18 18 46 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4455 $Y2=0.0360
r19 45 46 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4455 $Y2=0.0360
r20 44 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4185
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r21 43 44 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0360 $X2=0.4185 $Y2=0.0360
r22 42 43 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3800
+ $Y=0.0360 $X2=0.4050 $Y2=0.0360
r23 41 42 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3620
+ $Y=0.0360 $X2=0.3800 $Y2=0.0360
r24 40 41 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0360 $X2=0.3620 $Y2=0.0360
r25 39 40 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.0360 $X2=0.3510 $Y2=0.0360
r26 38 39 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.3240 $Y2=0.0360
r27 37 38 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2860
+ $Y=0.0360 $X2=0.2970 $Y2=0.0360
r28 36 37 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2680
+ $Y=0.0360 $X2=0.2860 $Y2=0.0360
r29 35 36 4.13912 $w=1.3e-08 $l=1.78e-08 $layer=M1 $thickness=3.6e-08 $X=0.2502
+ $Y=0.0360 $X2=0.2680 $Y2=0.0360
r30 34 35 0.524677 $w=1.3e-08 $l=2.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.2480
+ $Y=0.0360 $X2=0.2502 $Y2=0.0360
r31 34 33 1.69063 $w=1.3e-08 $l=7.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.2480
+ $Y=0.0360 $X2=0.2407 $Y2=0.0360
r32 32 33 5.77145 $w=1.3e-08 $l=2.47e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.2407 $Y2=0.0360
r33 31 32 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r34 30 31 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1755
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r35 29 30 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r36 15 29 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1500
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r37 11 1 0.958606 $w=2.2e-08 $l=2.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1640 $Y=0.0945 $X2=0.1640 $Y2=0.0725
r38 1 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r39 24 1 0.705882 $w=1.7e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1520 $Y=0.0725 $X2=0.1640 $Y2=0.0725
r40 13 24 0.264706 $w=1.7e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0725 $X2=0.1520 $Y2=0.0725
r41 13 1 0.471383 $w=3.35517e-08 $l=3.06472e-08 $layer=N_src_drn
+ $thickness=1e-09 $X=0.1475 $Y=0.0725 $X2=0.1620 $Y2=0.0455
r42 23 21 0.0675676 $w=3.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0455 $X2=0.1765 $Y2=0.0455
r43 1 21 0.391892 $w=3.7e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.0455 $X2=0.1765 $Y2=0.0455
r44 1 24 0.441971 $w=3.41429e-08 $l=2.87924e-08 $layer=N_src_drn
+ $thickness=1e-09 $X=0.1620 $Y=0.0455 $X2=0.1520 $Y2=0.0725
r45 10 1 0.391892 $w=3.7e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0455 $X2=0.1620 $Y2=0.0455
r46 22 10 0.0675676 $w=3.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0455 $X2=0.1475 $Y2=0.0455
r47 1 11 1e-05
.ends

.subckt PM_AOI322xp5_ASAP7_75t_R%NET53 VSS 16 17 31 34 36 10 1 11 2 12 3 13
c1 1 VSS 0.00458481f
c2 2 VSS 0.00461198f
c3 3 VSS 0.00507465f
c4 10 VSS 0.00216443f
c5 11 VSS 0.00216718f
c6 12 VSS 0.00221544f
c7 13 VSS 0.0214015f
r1 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4300 $Y2=0.2025
r2 36 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r3 34 33 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r4 32 33 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3340 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r5 2 32 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3220 $Y=0.2025 $X2=0.3340 $Y2=0.2025
r6 11 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3220 $Y2=0.2025
r7 31 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r8 3 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.2340
r9 2 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.2340
r10 27 28 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3935
+ $Y=0.2340 $X2=0.4320 $Y2=0.2340
r11 26 27 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3620
+ $Y=0.2340 $X2=0.3935 $Y2=0.2340
r12 25 26 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.2340 $X2=0.3620 $Y2=0.2340
r13 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.2340 $X2=0.3510 $Y2=0.2340
r14 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.2340 $X2=0.3375 $Y2=0.2340
r15 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3105
+ $Y=0.2340 $X2=0.3240 $Y2=0.2340
r16 21 22 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.2340 $X2=0.3105 $Y2=0.2340
r17 20 21 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2860
+ $Y=0.2340 $X2=0.2970 $Y2=0.2340
r18 19 20 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2545
+ $Y=0.2340 $X2=0.2860 $Y2=0.2340
r19 18 19 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2545 $Y2=0.2340
r20 13 18 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2045
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r21 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.2340
r22 16 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r23 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r24 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r25 17 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
.ends


*
.SUBCKT AOI322xp5_ASAP7_75t_R VSS VDD B2 B1 A1 A2 A3 C2 C1 Y
*
* VSS VSS
* VDD VDD
* B2 B2
* B1 B1
* A1 A1
* A2 A2
* A3 A3
* C2 C2
* C1 C1
* Y Y
*
*

MM4 N_MM4_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g N_MM3_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM0 N_MM0_d N_MM0_g N_MM0_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM11_g N_MM1_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM13_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM12_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM9_g N_MM5_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM10 N_MM10_d N_MM4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM0_g N_MM8_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 N_MM11_d N_MM11_g N_MM11_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM13 N_MM13_d N_MM13_g N_MM13_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM12 N_MM12_d N_MM12_g N_MM12_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g N_MM9_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AOI322xp5_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AOI322xp5_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AOI322xp5_ASAP7_75t_R%NET52 VSS N_MM1_s N_MM2_d N_NET52_1
+ PM_AOI322xp5_ASAP7_75t_R%NET52
cc_1 N_NET52_1 N_MM11_g 0.0173987f
cc_2 N_NET52_1 N_MM13_g 0.0172977f
x_PM_AOI322xp5_ASAP7_75t_R%NET51 VSS N_MM4_d N_MM3_s N_NET51_1
+ PM_AOI322xp5_ASAP7_75t_R%NET51
cc_3 N_NET51_1 N_MM4_g 0.0126231f
cc_4 N_NET51_1 N_MM3_g 0.0125589f
x_PM_AOI322xp5_ASAP7_75t_R%NET50 VSS N_MM6_d N_MM5_s N_NET50_1
+ PM_AOI322xp5_ASAP7_75t_R%NET50
cc_5 N_NET50_1 N_MM12_g 0.0126487f
cc_6 N_NET50_1 N_MM9_g 0.0125769f
x_PM_AOI322xp5_ASAP7_75t_R%NET49 VSS N_MM0_s N_MM1_d N_NET49_1
+ PM_AOI322xp5_ASAP7_75t_R%NET49
cc_7 N_NET49_1 N_MM0_g 0.0172956f
cc_8 N_NET49_1 N_MM11_g 0.0172811f
x_PM_AOI322xp5_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_AOI322xp5_ASAP7_75t_R%noxref_18
cc_9 N_noxref_18_1 N_MM4_g 0.00173505f
cc_10 N_noxref_18_1 N_NET27_10 0.0364059f
cc_11 N_noxref_18_1 N_noxref_17_1 0.00192f
x_PM_AOI322xp5_ASAP7_75t_R%B2 VSS B2 N_MM4_g N_B2_1 N_B2_4
+ PM_AOI322xp5_ASAP7_75t_R%B2
x_PM_AOI322xp5_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_AOI322xp5_ASAP7_75t_R%noxref_17
cc_12 N_noxref_17_1 N_MM4_g 0.00372059f
cc_13 N_noxref_17_1 N_NET27_10 0.000742177f
x_PM_AOI322xp5_ASAP7_75t_R%B1 VSS B1 N_MM3_g N_B1_1 N_B1_4
+ PM_AOI322xp5_ASAP7_75t_R%B1
cc_14 N_B1_1 N_B2_1 0.00134177f
cc_15 N_B1_4 N_B2_4 0.00402109f
cc_16 N_MM3_g N_MM4_g 0.00758512f
x_PM_AOI322xp5_ASAP7_75t_R%A3 VSS A3 N_MM13_g N_A3_1 N_A3_4
+ PM_AOI322xp5_ASAP7_75t_R%A3
cc_17 N_A3_1 N_A2_1 0.00129561f
cc_18 N_A3_4 N_A2_4 0.00336075f
cc_19 N_MM13_g N_MM11_g 0.00602807f
x_PM_AOI322xp5_ASAP7_75t_R%C2 VSS C2 N_MM12_g N_C2_4 N_C2_1
+ PM_AOI322xp5_ASAP7_75t_R%C2
cc_20 N_C2_4 N_A3_1 0.00085727f
cc_21 N_MM12_g N_MM13_g 0.00326931f
cc_22 N_C2_4 N_A3_4 0.00413983f
x_PM_AOI322xp5_ASAP7_75t_R%A2 VSS A2 N_MM11_g N_A2_1 N_A2_4
+ PM_AOI322xp5_ASAP7_75t_R%A2
cc_23 N_A2_1 N_A1_1 0.00122123f
cc_24 N_A2_4 N_A1_4 0.00343749f
cc_25 N_MM11_g N_MM0_g 0.00609968f
x_PM_AOI322xp5_ASAP7_75t_R%A1 VSS A1 N_MM0_g N_A1_1 N_A1_4
+ PM_AOI322xp5_ASAP7_75t_R%A1
cc_26 N_A1_1 N_MM3_g 0.000871754f
cc_27 N_A1_4 N_B1_4 0.00316964f
cc_28 N_MM0_g N_MM3_g 0.00399581f
x_PM_AOI322xp5_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_AOI322xp5_ASAP7_75t_R%noxref_19
cc_29 N_noxref_19_1 N_MM9_g 0.00350148f
cc_30 N_noxref_19_1 N_NET53_12 0.000584754f
cc_31 N_noxref_19_1 N_Y_12 0.0278821f
x_PM_AOI322xp5_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_AOI322xp5_ASAP7_75t_R%noxref_20
cc_32 N_noxref_20_1 N_MM9_g 0.00159439f
cc_33 N_noxref_20_1 N_NET53_12 0.036327f
cc_34 N_noxref_20_1 N_Y_14 0.00087312f
cc_35 N_noxref_20_1 N_noxref_19_1 0.00190183f
x_PM_AOI322xp5_ASAP7_75t_R%NET27 VSS N_MM11_s N_MM13_s N_MM7_d N_MM8_s N_MM10_d
+ N_NET27_10 N_NET27_1 N_NET27_13 N_NET27_11 N_NET27_2 N_NET27_12 N_NET27_3
+ PM_AOI322xp5_ASAP7_75t_R%NET27
cc_36 N_NET27_10 N_B2_1 0.000830406f
cc_37 N_NET27_1 N_MM4_g 0.00117899f
cc_38 N_NET27_13 N_B2_4 0.00147322f
cc_39 N_NET27_1 N_B2_4 0.0016648f
cc_40 N_NET27_10 N_MM4_g 0.0346438f
cc_41 N_NET27_11 N_B1_1 0.000798099f
cc_42 N_NET27_2 N_MM3_g 0.0008713f
cc_43 N_NET27_13 N_B1_4 0.00128908f
cc_44 N_NET27_2 N_B1_4 0.00131054f
cc_45 N_NET27_11 N_MM3_g 0.0339348f
cc_46 N_NET27_11 N_A1_1 0.000761917f
cc_47 N_NET27_2 N_MM0_g 0.00086441f
cc_48 N_NET27_13 N_A1_4 0.00125316f
cc_49 N_NET27_2 N_A1_4 0.00130046f
cc_50 N_NET27_11 N_MM0_g 0.0339987f
cc_51 N_NET27_12 N_A2_1 0.000680543f
cc_52 N_NET27_3 N_MM11_g 0.000888555f
cc_53 N_NET27_13 N_A2_4 0.00121151f
cc_54 N_NET27_3 N_A2_4 0.0012491f
cc_55 N_NET27_12 N_MM11_g 0.0340467f
cc_56 N_NET27_12 N_A3_4 0.000618488f
cc_57 N_NET27_12 N_A3_1 0.00076441f
cc_58 N_NET27_3 N_A3_4 0.00077809f
cc_59 N_NET27_3 N_MM13_g 0.000897818f
cc_60 N_NET27_12 N_MM13_g 0.0337883f
x_PM_AOI322xp5_ASAP7_75t_R%C1 VSS C1 N_MM9_g N_C1_1 N_C1_4
+ PM_AOI322xp5_ASAP7_75t_R%C1
cc_61 N_C1_1 N_C2_1 0.00120552f
cc_62 N_C1_4 N_C2_4 0.00334669f
cc_63 N_MM9_g N_MM12_g 0.00753327f
x_PM_AOI322xp5_ASAP7_75t_R%Y VSS Y N_MM3_d N_MM0_d N_MM5_d N_MM12_d N_MM9_d
+ N_Y_15 N_Y_10 N_Y_1 N_Y_11 N_Y_16 N_Y_14 N_Y_2 N_Y_3 N_Y_12 N_Y_17 N_Y_19
+ PM_AOI322xp5_ASAP7_75t_R%Y
cc_64 N_Y_15 N_MM3_g 0.000583331f
cc_65 N_Y_10 N_B1_1 0.000836265f
cc_66 N_Y_1 N_B1_4 0.00119382f
cc_67 N_Y_1 N_MM3_g 0.00155534f
cc_68 N_Y_11 N_MM3_g 0.00525961f
cc_69 N_Y_10 N_MM3_g 0.0303777f
cc_70 N_Y_10 N_A1_1 0.00066078f
cc_71 N_Y_15 N_A1_4 0.00126059f
cc_72 N_Y_1 N_MM0_g 0.0015373f
cc_73 N_Y_1 N_A1_4 0.00171966f
cc_74 N_Y_10 N_MM0_g 0.00980996f
cc_75 N_Y_11 N_MM0_g 0.0248666f
cc_76 N_Y_15 N_A2_4 0.00393971f
cc_77 N_Y_15 N_A3_4 0.00313793f
cc_78 N_Y_16 N_C2_4 0.00058278f
cc_79 N_Y_14 N_C2_1 0.000837671f
cc_80 N_Y_2 N_MM12_g 0.000914061f
cc_81 N_Y_15 N_C2_4 0.0013693f
cc_82 N_Y_2 N_C2_4 0.00210489f
cc_83 N_Y_14 N_MM12_g 0.0353363f
cc_84 N_Y_2 N_C1_1 0.000704076f
cc_85 N_Y_2 N_MM9_g 0.000896561f
cc_86 N_Y_3 N_MM9_g 0.000940566f
cc_87 N_Y_16 N_C1_4 0.0010967f
cc_88 N_Y_14 N_C1_1 0.00119307f
cc_89 N_Y_15 N_C1_4 0.00124309f
cc_90 N_Y_12 N_MM9_g 0.0109415f
cc_91 N_Y_17 N_C1_4 0.00675142f
cc_92 N_Y_14 N_MM9_g 0.0487961f
cc_93 N_Y_14 N_NET53_13 0.000563614f
cc_94 N_Y_16 N_NET53_3 0.000630619f
cc_95 N_Y_19 N_NET53_13 0.000666416f
cc_96 N_Y_14 N_NET53_12 0.000710851f
cc_97 N_Y_17 N_NET53_3 0.000717963f
cc_98 N_Y_2 N_NET53_13 0.000965777f
cc_99 N_Y_14 N_NET53_11 0.0011274f
cc_100 N_Y_2 N_NET53_3 0.0024233f
cc_101 N_Y_2 N_NET53_2 0.00416396f
cc_102 N_Y_16 N_NET53_13 0.00875836f
x_PM_AOI322xp5_ASAP7_75t_R%NET53 VSS N_MM11_d N_MM8_d N_MM13_d N_MM12_s N_MM9_s
+ N_NET53_10 N_NET53_1 N_NET53_11 N_NET53_2 N_NET53_12 N_NET53_3 N_NET53_13
+ PM_AOI322xp5_ASAP7_75t_R%NET53
cc_103 N_NET53_10 N_A1_1 0.00069598f
cc_104 N_NET53_1 N_MM0_g 0.000893769f
cc_105 N_NET53_10 N_MM0_g 0.0340091f
cc_106 N_NET53_10 N_A2_1 0.000653828f
cc_107 N_NET53_1 N_MM11_g 0.000891936f
cc_108 N_NET53_10 N_MM11_g 0.0341211f
cc_109 N_NET53_11 N_A3_4 0.000446093f
cc_110 N_NET53_11 N_A3_1 0.000733955f
cc_111 N_NET53_2 N_MM13_g 0.000939629f
cc_112 N_NET53_11 N_MM13_g 0.0341689f
cc_113 N_NET53_11 N_C2_1 0.000754934f
cc_114 N_NET53_2 N_MM12_g 0.000933777f
cc_115 N_NET53_11 N_MM12_g 0.0344399f
cc_116 N_NET53_12 N_C1_1 0.000724447f
cc_117 N_NET53_3 N_MM9_g 0.00105428f
cc_118 N_NET53_12 N_MM9_g 0.0347348f
cc_119 N_NET53_11 N_NET27_12 0.000559937f
cc_120 N_NET53_1 N_NET27_13 0.000756479f
cc_121 N_NET53_13 N_NET27_3 0.000757266f
cc_122 N_NET53_10 N_NET27_12 0.00112787f
cc_123 N_NET53_10 N_NET27_11 0.0011297f
cc_124 N_NET53_2 N_NET27_3 0.00134089f
cc_125 N_NET53_1 N_NET27_3 0.00281623f
cc_126 N_NET53_1 N_NET27_2 0.00433326f
cc_127 N_NET53_13 N_NET27_13 0.0102704f
*END of AOI322xp5_ASAP7_75t_R.pxi
.ENDS
** Design:	AOI32xp33_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AOI32xp33_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AOI32xp33_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AOI32xp33_ASAP7_75t_R%NET26 VSS 2 3 1
c1 1 VSS 0.000879816f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0540 $X2=0.2700 $Y2=0.0540
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0540 $X2=0.2700 $Y2=0.0540
.ends

.subckt PM_AOI32xp33_ASAP7_75t_R%NET24 VSS 2 3 1
c1 1 VSS 0.000925051f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_AOI32xp33_ASAP7_75t_R%NET25 VSS 2 3 1
c1 1 VSS 0.000900468f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_AOI32xp33_ASAP7_75t_R%B2 VSS 6 3 1 4
c1 1 VSS 0.00488467f
c2 3 VSS 0.00764674f
c3 4 VSS 0.00331772f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.0980
r2 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_AOI32xp33_ASAP7_75t_R%A1 VSS 23 3 9 7 6 1 4
c1 1 VSS 0.00178324f
c2 3 VSS 0.0327781f
c3 4 VSS 0.00324015f
c4 5 VSS 0.00768972f
c5 6 VSS 0.00172589f
c6 7 VSS 0.00286702f
c7 8 VSS 0.00175842f
c8 9 VSS 0.00812158f
r1 23 9 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0357
+ $Y=0.2340 $X2=0.0267 $Y2=0.2340
r2 23 20 2.12422 $w=1.31351e-08 $l=1.99922e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0357 $Y=0.2340 $X2=0.0270 $Y2=0.2160
r3 19 20 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1980 $X2=0.0270 $Y2=0.2160
r4 5 8 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1665 $X2=0.0270 $Y2=0.1350
r5 5 19 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1665 $X2=0.0270 $Y2=0.1980
r6 4 8 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1035 $X2=0.0270 $Y2=0.1350
r7 4 7 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1035 $X2=0.0270 $Y2=0.0720
r8 16 17 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0565
+ $Y=0.1350 $X2=0.0655 $Y2=0.1350
r9 6 16 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0455
+ $Y=0.1350 $X2=0.0565 $Y2=0.1350
r10 6 8 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0455 $Y=0.1350 $X2=0.0270 $Y2=0.1350
r11 14 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0605 $Y=0.1350
+ $X2=0.0655 $Y2=0.1350
r12 12 14 4.72579 $w=1.53e-08 $l=8e-09 $layer=LIG $thickness=4.8e-08 $X=0.0685
+ $Y=0.1350 $X2=0.0605 $Y2=0.1350
r13 1 11 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.0720
+ $Y=0.1350 $X2=0.0820 $Y2=0.1350
r14 1 12 1.73797 $w=1.72143e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0720 $Y=0.1350 $X2=0.0685 $Y2=0.1350
r15 3 11 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0820 $Y2=0.1350
r16 3 12 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0685 $Y2=0.1350
.ends

.subckt PM_AOI32xp33_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.0316193f
.ends

.subckt PM_AOI32xp33_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00452402f
.ends

.subckt PM_AOI32xp33_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.0048174f
.ends

.subckt PM_AOI32xp33_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.00500285f
.ends

.subckt PM_AOI32xp33_ASAP7_75t_R%A3 VSS 11 3 1 4 5
c1 1 VSS 0.00526829f
c2 3 VSS 0.0723437f
c3 4 VSS 0.00374097f
c4 5 VSS 0.00209642f
r1 11 5 0.382667 $w=1.8e-08 $l=3.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.1870
+ $Y=0.1980 $X2=0.1832 $Y2=0.1980
r2 11 10 2.96589 $w=1.31923e-08 $l=2.15928e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1870 $Y=0.1980 $X2=0.1890 $Y2=0.1765
r3 8 10 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1540 $X2=0.1890 $Y2=0.1765
r4 7 8 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1540
r5 4 7 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1035 $X2=0.1890 $Y2=0.1350
r6 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r7 1 7 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AOI32xp33_ASAP7_75t_R%B1 VSS 6 3 1 4
c1 1 VSS 0.00562755f
c2 3 VSS 0.0456326f
c3 4 VSS 0.00372636f
r1 7 8 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1230 $X2=0.2430 $Y2=0.1350
r2 6 7 0.816164 $w=1.3e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1195 $X2=0.2430 $Y2=0.1230
r3 6 4 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1195 $X2=0.2430 $Y2=0.0945
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AOI32xp33_ASAP7_75t_R%A2 VSS 10 3 1 6 5 4
c1 1 VSS 0.00337561f
c2 3 VSS 0.0349276f
c3 4 VSS 0.00256619f
c4 5 VSS 0.00205309f
c5 6 VSS 0.00228445f
r1 6 9 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1980 $X2=0.1350 $Y2=0.1665
r2 10 5 0.484711 $w=1.8e-08 $l=4.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0720 $X2=0.1302 $Y2=0.0720
r3 10 8 5.29779 $w=1.31087e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.0720 $X2=0.1350 $Y2=0.1035
r4 4 8 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1035
r5 4 9 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1665
r6 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r7 1 4 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AOI32xp33_ASAP7_75t_R%Y VSS 37 19 43 51 52 1 10 13 14 12 2 15 3 11 17
c1 1 VSS 0.00591551f
c2 2 VSS 0.0027756f
c3 3 VSS 0.00557636f
c4 10 VSS 0.00267847f
c5 11 VSS 0.002626f
c6 12 VSS 0.00215235f
c7 13 VSS 0.0285888f
c8 14 VSS 0.000657544f
c9 15 VSS 0.00208398f
c10 16 VSS 0.00282425f
c11 17 VSS 0.000768693f
r1 52 50 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2160 $X2=0.2845 $Y2=0.2160
r2 2 50 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.2160 $X2=0.2845 $Y2=0.2160
r3 12 2 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2160 $X2=0.2700 $Y2=0.2160
r4 51 12 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2160 $X2=0.2555 $Y2=0.2160
r5 2 47 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2160
+ $X2=0.2700 $Y2=0.1980
r6 47 48 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1980 $X2=0.2835 $Y2=0.1980
r7 45 48 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1980 $X2=0.2835 $Y2=0.1980
r8 44 45 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3220
+ $Y=0.1980 $X2=0.2970 $Y2=0.1980
r9 14 17 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3400 $Y=0.1980 $X2=0.3510 $Y2=0.1980
r10 14 44 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3400
+ $Y=0.1980 $X2=0.3220 $Y2=0.1980
r11 17 41 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.1980 $X2=0.3510 $Y2=0.1765
r12 11 3 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0540 $X2=0.3220 $Y2=0.0540
r13 43 11 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0540 $X2=0.3095 $Y2=0.0540
r14 40 41 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1170 $X2=0.3510 $Y2=0.1765
r15 39 40 11.7761 $w=1.3e-08 $l=5.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0665 $X2=0.3510 $Y2=0.1170
r16 15 38 2.63444 $w=1.48421e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.0540 $X2=0.3510 $Y2=0.0397
r17 15 39 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0540 $X2=0.3510 $Y2=0.0665
r18 3 35 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0540
+ $X2=0.3240 $Y2=0.0360
r19 37 38 0.586756 $w=1.8e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0340 $X2=0.3510 $Y2=0.0397
r20 37 16 0.382667 $w=1.8e-08 $l=3.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0340 $X2=0.3510 $Y2=0.0302
r21 37 36 1.10038 $w=5e-09 $l=1.36473e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.0340 $X2=0.3375 $Y2=0.0360
r22 35 36 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.0360 $X2=0.3375 $Y2=0.0360
r23 34 35 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3105
+ $Y=0.0360 $X2=0.3240 $Y2=0.0360
r24 33 34 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.3105 $Y2=0.0360
r25 32 33 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2720
+ $Y=0.0360 $X2=0.2970 $Y2=0.0360
r26 31 32 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2540
+ $Y=0.0360 $X2=0.2720 $Y2=0.0360
r27 30 31 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2540 $Y2=0.0360
r28 29 30 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2280
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r29 28 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2100
+ $Y=0.0360 $X2=0.2280 $Y2=0.0360
r30 27 28 4.89699 $w=1.3e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.2100 $Y2=0.0360
r31 26 27 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r32 25 26 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1240
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r33 24 25 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.0990
+ $Y=0.0360 $X2=0.1240 $Y2=0.0360
r34 23 24 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.0860
+ $Y=0.0360 $X2=0.0990 $Y2=0.0360
r35 22 23 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.0705
+ $Y=0.0360 $X2=0.0860 $Y2=0.0360
r36 21 22 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0605
+ $Y=0.0360 $X2=0.0705 $Y2=0.0360
r37 20 21 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0515
+ $Y=0.0360 $X2=0.0605 $Y2=0.0360
r38 13 20 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.0360 $X2=0.0515 $Y2=0.0360
r39 1 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0515 $Y2=0.0360
r40 19 18 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r41 10 18 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r42 1 10 1e-05
.ends

.subckt PM_AOI32xp33_ASAP7_75t_R%NET10 VSS 16 17 32 35 37 1 13 10 2 11 12 3
c1 1 VSS 0.00848586f
c2 2 VSS 0.00640677f
c3 3 VSS 0.00524263f
c4 10 VSS 0.00390045f
c5 11 VSS 0.00293844f
c6 12 VSS 0.0023317f
c7 13 VSS 0.0221755f
r1 12 3 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2160 $X2=0.3220 $Y2=0.2160
r2 37 12 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2160 $X2=0.3095 $Y2=0.2160
r3 35 34 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2160 $X2=0.2305 $Y2=0.2160
r4 33 34 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2260 $Y=0.2160 $X2=0.2305 $Y2=0.2160
r5 2 33 0.222222 $w=5.4e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2140 $Y=0.2160 $X2=0.2260 $Y2=0.2160
r6 11 2 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2160 $X2=0.2140 $Y2=0.2160
r7 32 11 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2160 $X2=0.2015 $Y2=0.2160
r8 3 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2160
+ $X2=0.3240 $Y2=0.2340
r9 2 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2160
+ $X2=0.2145 $Y2=0.2340
r10 28 29 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2855
+ $Y=0.2340 $X2=0.3240 $Y2=0.2340
r11 27 28 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2540
+ $Y=0.2340 $X2=0.2855 $Y2=0.2340
r12 26 27 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2540 $Y2=0.2340
r13 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.2340 $X2=0.2430 $Y2=0.2340
r14 24 25 1.39914 $w=1.3e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.2235
+ $Y=0.2340 $X2=0.2295 $Y2=0.2340
r15 23 24 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2145
+ $Y=0.2340 $X2=0.2235 $Y2=0.2340
r16 22 23 4.89699 $w=1.3e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1935
+ $Y=0.2340 $X2=0.2145 $Y2=0.2340
r17 21 22 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1935 $Y2=0.2340
r18 20 21 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1305
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r19 19 20 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1105
+ $Y=0.2340 $X2=0.1305 $Y2=0.2340
r20 18 19 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1015
+ $Y=0.2340 $X2=0.1105 $Y2=0.2340
r21 13 18 1.16595 $w=1.3e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0965
+ $Y=0.2340 $X2=0.1015 $Y2=0.2340
r22 1 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2160
+ $X2=0.1105 $Y2=0.2340
r23 17 15 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2160 $X2=0.1225 $Y2=0.2160
r24 1 15 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2160 $X2=0.1225 $Y2=0.2160
r25 10 1 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2160 $X2=0.1080 $Y2=0.2160
r26 16 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2160 $X2=0.0935 $Y2=0.2160
.ends


*
.SUBCKT AOI32xp33_ASAP7_75t_R VSS VDD A1 A2 A3 B1 B2 Y
*
* VSS VSS
* VDD VDD
* A1 A1
* A2 A2
* A3 A3
* B1 B1
* B2 B2
* Y Y
*
*

MM0 N_MM0_d N_MM0_g N_MM0_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM13 VSS N_MM13_g N_MM13_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM18 N_MM18_d N_MM18_g N_MM18_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1 N_MM1_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM4 N_MM4_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM14 N_MM14_d N_MM13_g N_MM14_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM15 N_MM15_d N_MM18_g N_MM15_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2


*include "AOI32xp33_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AOI32xp33_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AOI32xp33_ASAP7_75t_R%NET26 VSS N_MM13_s N_MM18_d N_NET26_1
+ PM_AOI32xp33_ASAP7_75t_R%NET26
cc_1 N_NET26_1 N_MM13_g 0.0125707f
cc_2 N_NET26_1 N_MM18_g 0.0125241f
x_PM_AOI32xp33_ASAP7_75t_R%NET24 VSS N_MM0_s N_MM2_d N_NET24_1
+ PM_AOI32xp33_ASAP7_75t_R%NET24
cc_3 N_NET24_1 N_MM0_g 0.0174552f
cc_4 N_NET24_1 N_MM2_g 0.0174156f
x_PM_AOI32xp33_ASAP7_75t_R%NET25 VSS N_MM2_s N_MM3_d N_NET25_1
+ PM_AOI32xp33_ASAP7_75t_R%NET25
cc_5 N_NET25_1 N_MM2_g 0.0174536f
cc_6 N_NET25_1 N_MM3_g 0.0173419f
x_PM_AOI32xp33_ASAP7_75t_R%B2 VSS B2 N_MM18_g N_B2_1 N_B2_4
+ PM_AOI32xp33_ASAP7_75t_R%B2
cc_7 N_B2_1 N_B1_1 0.00162993f
cc_8 N_B2_4 N_B1_4 0.00368415f
cc_9 N_MM18_g N_MM13_g 0.00968945f
x_PM_AOI32xp33_ASAP7_75t_R%A1 VSS A1 N_MM0_g N_A1_9 N_A1_7 N_A1_6 N_A1_1 N_A1_4
+ PM_AOI32xp33_ASAP7_75t_R%A1
x_PM_AOI32xp33_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_AOI32xp33_ASAP7_75t_R%noxref_14
cc_10 N_noxref_14_1 N_MM0_g 0.00469448f
cc_11 N_noxref_14_1 N_Y_10 0.000494292f
cc_12 N_noxref_14_1 N_noxref_13_1 0.00185822f
x_PM_AOI32xp33_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_AOI32xp33_ASAP7_75t_R%noxref_15
cc_13 N_noxref_15_1 N_MM18_g 0.00368749f
cc_14 N_noxref_15_1 N_Y_11 0.0283482f
x_PM_AOI32xp33_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_AOI32xp33_ASAP7_75t_R%noxref_13
cc_15 N_noxref_13_1 N_MM0_g 0.0025574f
cc_16 N_noxref_13_1 N_Y_10 0.0371547f
x_PM_AOI32xp33_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_AOI32xp33_ASAP7_75t_R%noxref_16
cc_17 N_noxref_16_1 N_MM18_g 0.00366441f
cc_18 N_noxref_16_1 N_NET10_12 0.0267692f
cc_19 N_noxref_16_1 N_Y_12 0.00109231f
cc_20 N_noxref_16_1 N_noxref_15_1 0.00205173f
x_PM_AOI32xp33_ASAP7_75t_R%A3 VSS A3 N_MM3_g N_A3_1 N_A3_4 N_A3_5
+ PM_AOI32xp33_ASAP7_75t_R%A3
cc_21 N_MM3_g N_A2_6 0.000874488f
cc_22 N_A3_1 N_A2_1 0.0027972f
cc_23 N_A3_4 N_A2_4 0.0043585f
cc_24 N_MM3_g N_MM2_g 0.00762878f
x_PM_AOI32xp33_ASAP7_75t_R%B1 VSS B1 N_MM13_g N_B1_1 N_B1_4
+ PM_AOI32xp33_ASAP7_75t_R%B1
cc_25 N_B1_1 N_A3_1 0.001258f
cc_26 N_B1_4 N_A3_4 0.0039927f
cc_27 N_MM13_g N_MM3_g 0.0066429f
x_PM_AOI32xp33_ASAP7_75t_R%A2 VSS A2 N_MM2_g N_A2_1 N_A2_6 N_A2_5 N_A2_4
+ PM_AOI32xp33_ASAP7_75t_R%A2
cc_28 N_A2_1 N_MM0_g 0.000394923f
cc_29 N_A2_6 N_A1_9 0.000638568f
cc_30 N_A2_5 N_A1_7 0.000825208f
cc_31 N_A2_4 N_A1_6 0.0018342f
cc_32 N_A2_1 N_A1_1 0.00188197f
cc_33 N_MM2_g N_MM0_g 0.00809372f
x_PM_AOI32xp33_ASAP7_75t_R%Y VSS Y N_MM0_d N_MM18_s N_MM14_d N_MM15_d N_Y_1
+ N_Y_10 N_Y_13 N_Y_14 N_Y_12 N_Y_2 N_Y_15 N_Y_3 N_Y_11 N_Y_17
+ PM_AOI32xp33_ASAP7_75t_R%Y
cc_34 N_Y_1 N_MM0_g 0.00310383f
cc_35 N_Y_1 N_A1_4 0.00051233f
cc_36 N_Y_10 N_A1_1 0.00179302f
cc_37 N_Y_13 N_A1_7 0.00370882f
cc_38 N_Y_10 N_MM0_g 0.0366243f
cc_39 N_Y_1 N_A2_5 0.000434127f
cc_40 N_Y_13 N_A2_4 0.000449089f
cc_41 N_Y_13 N_A2_5 0.00627923f
cc_42 N_Y_14 N_A3_4 0.000775098f
cc_43 N_Y_13 N_A3_4 0.00321721f
cc_44 N_Y_12 N_B1_1 0.000349679f
cc_45 N_Y_2 N_MM13_g 0.000463371f
cc_46 N_Y_14 N_B1_4 0.000570674f
cc_47 N_Y_13 N_B1_4 0.00349255f
cc_48 N_Y_12 N_MM13_g 0.0261585f
cc_49 N_Y_2 N_MM18_g 0.000458374f
cc_50 N_Y_15 N_B2_1 0.000641196f
cc_51 N_Y_12 N_B2_1 0.000853354f
cc_52 N_Y_3 N_MM18_g 0.000960742f
cc_53 N_Y_14 N_B2_4 0.00120355f
cc_54 N_Y_13 N_B2_4 0.00122493f
cc_55 N_Y_12 N_MM18_g 0.01094f
cc_56 N_Y_15 N_B2_4 0.00669947f
cc_57 N_Y_11 N_MM18_g 0.0401101f
cc_58 N_Y_15 N_NET10_13 0.000471144f
cc_59 N_Y_12 N_NET10_12 0.000524044f
cc_60 N_Y_17 N_NET10_13 0.000578743f
cc_61 N_Y_2 N_NET10_13 0.000653026f
cc_62 N_Y_14 N_NET10_3 0.000668809f
cc_63 N_Y_12 N_NET10_11 0.00083162f
cc_64 N_Y_2 N_NET10_3 0.00171041f
cc_65 N_Y_2 N_NET10_2 0.00304279f
cc_66 N_Y_14 N_NET10_13 0.00857145f
x_PM_AOI32xp33_ASAP7_75t_R%NET10 VSS N_MM5_d N_MM1_d N_MM4_d N_MM14_s N_MM15_s
+ N_NET10_1 N_NET10_13 N_NET10_10 N_NET10_2 N_NET10_11 N_NET10_12 N_NET10_3
+ PM_AOI32xp33_ASAP7_75t_R%NET10
cc_67 N_NET10_1 N_MM0_g 0.000581538f
cc_68 N_NET10_13 N_A1_9 0.000913522f
cc_69 N_NET10_10 N_MM0_g 0.0252761f
cc_70 N_NET10_10 N_A2_4 0.000426437f
cc_71 N_NET10_1 N_MM2_g 0.000859875f
cc_72 N_NET10_13 N_A2_6 0.00448969f
cc_73 N_NET10_10 N_MM2_g 0.0250608f
cc_74 N_NET10_2 N_MM3_g 0.000807466f
cc_75 N_NET10_13 N_A3_5 0.00492784f
cc_76 N_NET10_11 N_MM3_g 0.0255725f
cc_77 N_NET10_11 N_MM13_g 0.025558f
cc_78 N_NET10_12 N_MM18_g 0.0256104f
*END of AOI32xp33_ASAP7_75t_R.pxi
.ENDS
** Design:	AOI331xp33_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AOI331xp33_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AOI331xp33_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AOI331xp33_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.0429086f
.ends

.subckt PM_AOI331xp33_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.042835f
.ends

.subckt PM_AOI331xp33_ASAP7_75t_R%NET25 VSS 2 3 1
c1 1 VSS 0.000950527f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_AOI331xp33_ASAP7_75t_R%NET064 VSS 2 3 1
c1 1 VSS 0.000960013f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3240 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3240 $Y2=0.0675
.ends

.subckt PM_AOI331xp33_ASAP7_75t_R%NET063 VSS 2 3 1
c1 1 VSS 0.000994783f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2700 $Y2=0.0675
.ends

.subckt PM_AOI331xp33_ASAP7_75t_R%NET26 VSS 2 3 1
c1 1 VSS 0.000952716f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_AOI331xp33_ASAP7_75t_R%A3 VSS 6 3 1 4
c1 1 VSS 0.00557185f
c2 3 VSS 0.0821009f
c3 4 VSS 0.0187108f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1207 $X2=0.0810 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1150 $X2=0.0810 $Y2=0.1207
r3 6 4 9.50248 $w=1.3e-08 $l=4.08e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1150 $X2=0.0810 $Y2=0.0742
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AOI331xp33_ASAP7_75t_R%A2 VSS 6 3 1 4
c1 1 VSS 0.00681621f
c2 3 VSS 0.0472754f
c3 4 VSS 0.00900259f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1207 $X2=0.1350 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1150 $X2=0.1350 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1150 $X2=0.1350 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AOI331xp33_ASAP7_75t_R%NET031 VSS 16 17 34 35 38 39 10 1 13 2 11 12 3
c1 1 VSS 0.00999362f
c2 2 VSS 0.00695531f
c3 3 VSS 0.00458308f
c4 10 VSS 0.00461067f
c5 11 VSS 0.00338049f
c6 12 VSS 0.00217925f
c7 13 VSS 0.0217928f
r1 39 37 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r2 3 37 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r3 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r4 38 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r5 35 33 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r6 1 33 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r7 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r8 34 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
r9 3 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.2340
r10 1 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.2340
r11 29 30 9.211 $w=1.3e-08 $l=3.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2845
+ $Y=0.2340 $X2=0.3240 $Y2=0.2340
r12 28 29 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2530
+ $Y=0.2340 $X2=0.2845 $Y2=0.2340
r13 27 28 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2530 $Y2=0.2340
r14 26 27 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.2340 $X2=0.2430 $Y2=0.2340
r15 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2295 $Y2=0.2340
r16 24 25 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2040
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r17 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.1215 $Y2=0.2340
r18 20 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1215 $Y2=0.2340
r19 19 20 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r20 18 19 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r21 13 18 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1995
+ $Y=0.2340 $X2=0.1890 $Y2=0.2340
r22 13 24 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1995
+ $Y=0.2340 $X2=0.2040 $Y2=0.2340
r23 2 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.2340
r24 16 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r25 2 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r26 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r27 17 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
.ends

.subckt PM_AOI331xp33_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.00495929f
.ends

.subckt PM_AOI331xp33_ASAP7_75t_R%B3 VSS 6 3 1 4
c1 1 VSS 0.00798966f
c2 3 VSS 0.0468352f
c3 4 VSS 0.0050268f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1207 $X2=0.3510 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1150 $X2=0.3510 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1150 $X2=0.3510 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
.ends

.subckt PM_AOI331xp33_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.005072f
.ends

.subckt PM_AOI331xp33_ASAP7_75t_R%A1 VSS 6 3 1 4
c1 1 VSS 0.00802022f
c2 3 VSS 0.0461061f
c3 4 VSS 0.00595019f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1207 $X2=0.1890 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1150 $X2=0.1890 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1150 $X2=0.1890 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AOI331xp33_ASAP7_75t_R%C1 VSS 6 3 4 1
c1 1 VSS 0.00861678f
c2 3 VSS 0.0456442f
c3 4 VSS 0.00515389f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1207 $X2=0.4050 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1150 $X2=0.4050 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1150 $X2=0.4050 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
.ends

.subckt PM_AOI331xp33_ASAP7_75t_R%B2 VSS 6 3 1 4
c1 1 VSS 0.00766331f
c2 3 VSS 0.0100186f
c3 4 VSS 0.00501254f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1207 $X2=0.2970 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1150 $X2=0.2970 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1150 $X2=0.2970 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_AOI331xp33_ASAP7_75t_R%NET030 VSS 12 13 25 26 7 1 9 8 2
c1 1 VSS 0.00288033f
c2 2 VSS 0.00319071f
c3 7 VSS 0.00211725f
c4 8 VSS 0.00217625f
c5 9 VSS 0.00218116f
r1 26 24 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r2 2 24 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3780 $Y2=0.2025
r4 25 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r5 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.1980
r6 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3645
+ $Y=0.1980 $X2=0.3780 $Y2=0.1980
r7 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1980 $X2=0.3645 $Y2=0.1980
r8 18 19 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.3405
+ $Y=0.1980 $X2=0.3510 $Y2=0.1980
r9 17 18 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3225
+ $Y=0.1980 $X2=0.3405 $Y2=0.1980
r10 16 17 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1980 $X2=0.3225 $Y2=0.1980
r11 15 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2835
+ $Y=0.1980 $X2=0.2970 $Y2=0.1980
r12 14 15 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1980 $X2=0.2835 $Y2=0.1980
r13 9 14 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2575
+ $Y=0.1980 $X2=0.2700 $Y2=0.1980
r14 1 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.1980
r15 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r16 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r17 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r18 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
.ends

.subckt PM_AOI331xp33_ASAP7_75t_R%B1 VSS 6 3 1 4
c1 1 VSS 0.00821692f
c2 3 VSS 0.00939605f
c3 4 VSS 0.00523096f
r1 7 8 3.20636 $w=1.3e-08 $l=1.38e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1212 $X2=0.2430 $Y2=0.1350
r2 6 7 1.22425 $w=1.3e-08 $l=5.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1160 $X2=0.2430 $Y2=0.1212
r3 6 4 5.42166 $w=1.3e-08 $l=2.33e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1160 $X2=0.2430 $Y2=0.0927
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AOI331xp33_ASAP7_75t_R%Y VSS 37 19 20 43 48 13 10 1 2 3 12 14 11 15
c1 1 VSS 0.00708403f
c2 2 VSS 0.00743213f
c3 3 VSS 0.00538818f
c4 10 VSS 0.00343814f
c5 11 VSS 0.00352954f
c6 12 VSS 0.00232237f
c7 13 VSS 0.0242361f
c8 14 VSS 0.00292224f
c9 15 VSS 0.00569031f
c10 16 VSS 0.00280667f
r1 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4300 $Y2=0.2025
r2 48 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r3 3 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.2340
r4 45 46 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4455 $Y2=0.2340
r5 15 41 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4590 $Y2=0.2160
r6 15 46 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.2340 $X2=0.4455 $Y2=0.2340
r7 11 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0675 $X2=0.4300 $Y2=0.0675
r8 43 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4175 $Y2=0.0675
r9 40 41 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1980 $X2=0.4590 $Y2=0.2160
r10 39 40 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1765 $X2=0.4590 $Y2=0.1980
r11 38 39 7.17059 $w=1.3e-08 $l=3.08e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1457 $X2=0.4590 $Y2=0.1765
r12 37 38 4.37231 $w=1.3e-08 $l=1.87e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1270 $X2=0.4590 $Y2=0.1457
r13 37 36 6.70421 $w=1.3e-08 $l=2.88e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1270 $X2=0.4590 $Y2=0.0982
r14 14 16 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0575 $X2=0.4590 $Y2=0.0360
r15 14 36 9.50248 $w=1.3e-08 $l=4.07e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0575 $X2=0.4590 $Y2=0.0982
r16 2 34 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4320 $Y2=0.0360
r17 16 35 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4455 $Y2=0.0360
r18 34 35 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4455 $Y2=0.0360
r19 33 34 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4200
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r20 32 33 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4155
+ $Y=0.0360 $X2=0.4200 $Y2=0.0360
r21 31 32 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0360 $X2=0.4155 $Y2=0.0360
r22 30 31 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.3945
+ $Y=0.0360 $X2=0.4050 $Y2=0.0360
r23 29 30 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3765
+ $Y=0.0360 $X2=0.3945 $Y2=0.0360
r24 28 29 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0360 $X2=0.3765 $Y2=0.0360
r25 27 28 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.0360 $X2=0.3510 $Y2=0.0360
r26 26 27 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.3240 $Y2=0.0360
r27 25 26 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2710
+ $Y=0.0360 $X2=0.2970 $Y2=0.0360
r28 24 25 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2530
+ $Y=0.0360 $X2=0.2710 $Y2=0.0360
r29 23 24 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2530 $Y2=0.0360
r30 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r31 21 22 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.2295 $Y2=0.0360
r32 13 21 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2040
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r33 1 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0675
+ $X2=0.2160 $Y2=0.0360
r34 20 18 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r35 1 18 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r36 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r37 19 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2015 $Y2=0.0675
.ends


*
.SUBCKT AOI331xp33_ASAP7_75t_R VSS VDD A3 A2 A1 B1 B2 B3 C1 Y
*
* VSS VSS
* VDD VDD
* A3 A3
* A2 A2
* A1 A1
* B1 B1
* B2 B2
* B3 B3
* C1 C1
* Y Y
*
*

MM3 N_MM3_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM14 N_MM14_d N_MM14_g N_MM14_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM12 N_MM12_d N_MM6_g N_MM12_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 N_MM11_d N_MM5_g N_MM11_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM17 N_MM17_d N_MM1_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM14_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM6_g N_MM6_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g N_MM4_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AOI331xp33_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AOI331xp33_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AOI331xp33_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_AOI331xp33_ASAP7_75t_R%noxref_18
cc_1 N_noxref_18_1 N_MM3_g 0.00166218f
cc_2 N_noxref_18_1 N_noxref_17_1 0.00179371f
x_PM_AOI331xp33_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_AOI331xp33_ASAP7_75t_R%noxref_17
cc_3 N_noxref_17_1 N_MM3_g 0.00167963f
x_PM_AOI331xp33_ASAP7_75t_R%NET25 VSS N_MM3_d N_MM2_s N_NET25_1
+ PM_AOI331xp33_ASAP7_75t_R%NET25
cc_4 N_NET25_1 N_MM3_g 0.0173555f
cc_5 N_NET25_1 N_MM2_g 0.0172619f
x_PM_AOI331xp33_ASAP7_75t_R%NET064 VSS N_MM11_s N_MM10_d N_NET064_1
+ PM_AOI331xp33_ASAP7_75t_R%NET064
cc_6 N_NET064_1 N_MM5_g 0.0174027f
cc_7 N_NET064_1 N_MM4_g 0.0173094f
x_PM_AOI331xp33_ASAP7_75t_R%NET063 VSS N_MM12_s N_MM11_d N_NET063_1
+ PM_AOI331xp33_ASAP7_75t_R%NET063
cc_8 N_NET063_1 N_MM6_g 0.0173153f
cc_9 N_NET063_1 N_MM5_g 0.0172504f
x_PM_AOI331xp33_ASAP7_75t_R%NET26 VSS N_MM2_d N_MM14_s N_NET26_1
+ PM_AOI331xp33_ASAP7_75t_R%NET26
cc_10 N_NET26_1 N_MM2_g 0.0172815f
cc_11 N_NET26_1 N_MM14_g 0.0171674f
x_PM_AOI331xp33_ASAP7_75t_R%A3 VSS A3 N_MM3_g N_A3_1 N_A3_4
+ PM_AOI331xp33_ASAP7_75t_R%A3
x_PM_AOI331xp33_ASAP7_75t_R%A2 VSS A2 N_MM2_g N_A2_1 N_A2_4
+ PM_AOI331xp33_ASAP7_75t_R%A2
cc_12 N_A2_1 N_A3_1 0.00136193f
cc_13 N_MM2_g N_MM3_g 0.00524155f
cc_14 N_A2_4 N_A3_4 0.00762236f
x_PM_AOI331xp33_ASAP7_75t_R%NET031 VSS N_MM6_s N_MM9_d N_MM7_d N_MM8_d N_MM5_s
+ N_MM4_s N_NET031_10 N_NET031_1 N_NET031_13 N_NET031_2 N_NET031_11 N_NET031_12
+ N_NET031_3 PM_AOI331xp33_ASAP7_75t_R%NET031
cc_15 N_NET031_10 N_A3_1 0.000659424f
cc_16 N_NET031_1 N_MM3_g 0.00118245f
cc_17 N_NET031_1 N_A3_4 0.00119656f
cc_18 N_NET031_10 N_MM3_g 0.0342269f
cc_19 N_NET031_13 N_A2_4 0.00111437f
cc_20 N_NET031_1 N_MM2_g 0.00115671f
cc_21 N_NET031_1 N_A2_4 0.00154452f
cc_22 N_NET031_10 N_MM2_g 0.0343134f
cc_23 N_NET031_13 N_A1_4 0.00118386f
cc_24 N_NET031_2 N_MM14_g 0.00119207f
cc_25 N_NET031_2 N_A1_4 0.00173747f
cc_26 N_NET031_11 N_MM14_g 0.034359f
cc_27 N_NET031_11 N_B1_1 0.000731887f
cc_28 N_NET031_2 N_MM6_g 0.000941691f
cc_29 N_NET031_11 N_MM6_g 0.0339239f
cc_30 N_NET031_12 N_B2_1 0.000734669f
cc_31 N_NET031_3 N_MM5_g 0.000917452f
cc_32 N_NET031_12 N_MM5_g 0.0338048f
cc_33 N_NET031_12 N_B3_1 0.00069552f
cc_34 N_NET031_3 N_MM4_g 0.000907516f
cc_35 N_NET031_12 N_MM4_g 0.0335736f
x_PM_AOI331xp33_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_AOI331xp33_ASAP7_75t_R%noxref_19
cc_36 N_noxref_19_1 N_MM1_g 0.0014511f
cc_37 N_noxref_19_1 N_Y_11 0.03822f
x_PM_AOI331xp33_ASAP7_75t_R%B3 VSS B3 N_MM4_g N_B3_1 N_B3_4
+ PM_AOI331xp33_ASAP7_75t_R%B3
cc_38 N_B3_1 N_B2_1 0.00123273f
cc_39 N_B3_4 N_B2_4 0.00360336f
cc_40 N_MM4_g N_MM5_g 0.00610958f
x_PM_AOI331xp33_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_AOI331xp33_ASAP7_75t_R%noxref_20
cc_41 N_noxref_20_1 N_MM1_g 0.0014549f
cc_42 N_noxref_20_1 N_Y_12 0.0381211f
cc_43 N_noxref_20_1 N_noxref_19_1 0.00177438f
x_PM_AOI331xp33_ASAP7_75t_R%A1 VSS A1 N_MM14_g N_A1_1 N_A1_4
+ PM_AOI331xp33_ASAP7_75t_R%A1
cc_44 N_A1_1 N_A2_1 0.00139308f
cc_45 N_MM14_g N_MM2_g 0.0051796f
cc_46 N_A1_4 N_A2_4 0.0061902f
x_PM_AOI331xp33_ASAP7_75t_R%C1 VSS C1 N_MM1_g N_C1_4 N_C1_1
+ PM_AOI331xp33_ASAP7_75t_R%C1
cc_47 N_MM1_g N_B3_1 0.00082186f
cc_48 N_C1_4 N_B3_4 0.00329239f
cc_49 N_MM1_g N_MM4_g 0.00410965f
x_PM_AOI331xp33_ASAP7_75t_R%B2 VSS B2 N_MM5_g N_B2_1 N_B2_4
+ PM_AOI331xp33_ASAP7_75t_R%B2
cc_50 N_B2_1 N_B1_1 0.00132305f
cc_51 N_B2_4 N_B1_4 0.00340282f
cc_52 N_MM5_g N_MM6_g 0.00600832f
x_PM_AOI331xp33_ASAP7_75t_R%NET030 VSS N_MM6_d N_MM5_d N_MM4_d N_MM1_s
+ N_NET030_7 N_NET030_1 N_NET030_9 N_NET030_8 N_NET030_2
+ PM_AOI331xp33_ASAP7_75t_R%NET030
cc_53 N_NET030_7 N_B1_4 0.000620925f
cc_54 N_NET030_1 N_B1_4 0.00073821f
cc_55 N_NET030_7 N_B1_1 0.000741041f
cc_56 N_NET030_1 N_MM6_g 0.000880359f
cc_57 N_NET030_7 N_MM6_g 0.0332658f
cc_58 N_NET030_7 N_B2_1 0.000829119f
cc_59 N_NET030_1 N_MM5_g 0.00086926f
cc_60 N_NET030_9 N_B2_4 0.00110006f
cc_61 N_NET030_1 N_B2_4 0.00125065f
cc_62 N_NET030_7 N_MM5_g 0.0333091f
cc_63 N_NET030_8 N_B3_1 0.000734667f
cc_64 N_NET030_2 N_MM4_g 0.000866472f
cc_65 N_NET030_9 N_B3_4 0.00110879f
cc_66 N_NET030_2 N_B3_4 0.00120758f
cc_67 N_NET030_8 N_MM4_g 0.0334137f
cc_68 N_NET030_8 N_C1_1 0.000666545f
cc_69 N_NET030_2 N_C1_4 0.000781816f
cc_70 N_NET030_2 N_MM1_g 0.000878142f
cc_71 N_NET030_8 N_MM1_g 0.0338515f
cc_72 N_NET030_7 N_NET031_13 0.000551583f
cc_73 N_NET030_1 N_NET031_13 0.000697901f
cc_74 N_NET030_9 N_NET031_3 0.000794598f
cc_75 N_NET030_7 N_NET031_11 0.00110844f
cc_76 N_NET030_7 N_NET031_12 0.00110985f
cc_77 N_NET030_2 N_NET031_3 0.00122385f
cc_78 N_NET030_1 N_NET031_3 0.00299156f
cc_79 N_NET030_1 N_NET031_2 0.00407851f
cc_80 N_NET030_9 N_NET031_13 0.00973923f
x_PM_AOI331xp33_ASAP7_75t_R%B1 VSS B1 N_MM6_g N_B1_1 N_B1_4
+ PM_AOI331xp33_ASAP7_75t_R%B1
cc_81 N_B1_1 N_A1_4 0.000919735f
cc_82 N_MM6_g N_MM14_g 0.00327403f
cc_83 N_B1_4 N_A1_4 0.00450351f
x_PM_AOI331xp33_ASAP7_75t_R%Y VSS Y N_MM14_d N_MM12_d N_MM17_d N_MM1_d N_Y_13
+ N_Y_10 N_Y_1 N_Y_2 N_Y_3 N_Y_12 N_Y_14 N_Y_11 N_Y_15
+ PM_AOI331xp33_ASAP7_75t_R%Y
cc_84 N_Y_13 N_MM14_g 0.000603211f
cc_85 N_Y_10 N_A1_1 0.000940684f
cc_86 N_Y_1 N_A1_4 0.00125133f
cc_87 N_Y_1 N_MM14_g 0.00155718f
cc_88 N_Y_10 N_MM14_g 0.0353551f
cc_89 N_Y_10 N_B1_1 0.000785192f
cc_90 N_Y_13 N_B1_4 0.00123491f
cc_91 N_Y_1 N_MM6_g 0.00153406f
cc_92 N_Y_1 N_B1_4 0.00174289f
cc_93 N_Y_10 N_MM6_g 0.0353058f
cc_94 N_Y_13 N_B2_4 0.0039741f
cc_95 N_Y_13 N_B3_4 0.00323257f
cc_96 N_Y_2 N_C1_1 0.000835893f
cc_97 N_Y_3 N_MM1_g 0.00109638f
cc_98 N_Y_13 N_C1_4 0.00111833f
cc_99 N_Y_2 N_MM1_g 0.00132126f
cc_100 N_Y_12 N_C1_1 0.00162745f
cc_101 N_Y_12 N_MM1_g 0.0151178f
cc_102 N_Y_14 N_C1_4 0.00612753f
cc_103 N_Y_11 N_MM1_g 0.0542649f
cc_104 N_Y_12 N_NET030_8 0.00110499f
cc_105 N_Y_15 N_NET030_9 0.00122042f
cc_106 N_Y_3 N_NET030_2 0.00384101f
*END of AOI331xp33_ASAP7_75t_R.pxi
.ENDS
** Design:	AOI332xp33_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AOI332xp33_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AOI332xp33_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AOI332xp33_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.0429004f
.ends

.subckt PM_AOI332xp33_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.0429128f
.ends

.subckt PM_AOI332xp33_ASAP7_75t_R%NET061 VSS 2 3 1
c1 1 VSS 0.00101423f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4320 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4320 $Y2=0.0675
.ends

.subckt PM_AOI332xp33_ASAP7_75t_R%NET064 VSS 2 3 1
c1 1 VSS 0.000993108f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3240 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3240 $Y2=0.0675
.ends

.subckt PM_AOI332xp33_ASAP7_75t_R%NET063 VSS 2 3 1
c1 1 VSS 0.00101118f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2700 $Y2=0.0675
.ends

.subckt PM_AOI332xp33_ASAP7_75t_R%NET25 VSS 2 3 1
c1 1 VSS 0.000947137f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_AOI332xp33_ASAP7_75t_R%NET26 VSS 2 3 1
c1 1 VSS 0.0009487f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_AOI332xp33_ASAP7_75t_R%A2 VSS 6 3 1 4
c1 1 VSS 0.00688628f
c2 3 VSS 0.0472887f
c3 4 VSS 0.00811941f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1207 $X2=0.1350 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1150 $X2=0.1350 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1150 $X2=0.1350 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AOI332xp33_ASAP7_75t_R%A3 VSS 6 3 1 4
c1 1 VSS 0.00557691f
c2 3 VSS 0.0820907f
c3 4 VSS 0.0170248f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1207 $X2=0.0810 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1150 $X2=0.0810 $Y2=0.1207
r3 6 4 9.50248 $w=1.3e-08 $l=4.08e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1150 $X2=0.0810 $Y2=0.0742
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AOI332xp33_ASAP7_75t_R%NET031 VSS 16 17 36 37 40 41 13 1 10 2 11 12 3
c1 1 VSS 0.0087652f
c2 2 VSS 0.00591119f
c3 3 VSS 0.00304125f
c4 10 VSS 0.00452419f
c5 11 VSS 0.0033356f
c6 12 VSS 0.00212992f
c7 13 VSS 0.00786396f
r1 41 39 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r2 3 39 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r3 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r4 40 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r5 37 35 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r6 1 35 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r7 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r8 36 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
r9 3 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.1980
r10 1 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.1980
r11 31 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3105
+ $Y=0.1980 $X2=0.3240 $Y2=0.1980
r12 30 31 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1980 $X2=0.3105 $Y2=0.1980
r13 29 30 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2710
+ $Y=0.1980 $X2=0.2970 $Y2=0.1980
r14 28 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2530
+ $Y=0.1980 $X2=0.2710 $Y2=0.1980
r15 27 28 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1980 $X2=0.2530 $Y2=0.1980
r16 26 27 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.1980 $X2=0.2430 $Y2=0.1980
r17 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1980 $X2=0.2295 $Y2=0.1980
r18 24 25 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2040
+ $Y=0.1980 $X2=0.2160 $Y2=0.1980
r19 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.1980 $X2=0.1215 $Y2=0.1980
r20 20 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1980 $X2=0.1215 $Y2=0.1980
r21 19 20 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.1980 $X2=0.1350 $Y2=0.1980
r22 18 19 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1980 $X2=0.1620 $Y2=0.1980
r23 13 18 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1995
+ $Y=0.1980 $X2=0.1890 $Y2=0.1980
r24 13 24 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1995
+ $Y=0.1980 $X2=0.2040 $Y2=0.1980
r25 2 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.1980
r26 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r27 2 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r28 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r29 16 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
.ends

.subckt PM_AOI332xp33_ASAP7_75t_R%B2 VSS 6 3 1 4
c1 1 VSS 0.00727386f
c2 3 VSS 0.00976358f
c3 4 VSS 0.00482539f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1207 $X2=0.2970 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1150 $X2=0.2970 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1150 $X2=0.2970 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_AOI332xp33_ASAP7_75t_R%C1 VSS 6 3 1 4
c1 1 VSS 0.00783439f
c2 3 VSS 0.00908318f
c3 4 VSS 0.00481892f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1207 $X2=0.4590 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1150 $X2=0.4590 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1150 $X2=0.4590 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1350
+ $X2=0.4590 $Y2=0.1350
.ends

.subckt PM_AOI332xp33_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.00550024f
.ends

.subckt PM_AOI332xp33_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.00601767f
.ends

.subckt PM_AOI332xp33_ASAP7_75t_R%A1 VSS 6 3 1 4
c1 1 VSS 0.00788632f
c2 3 VSS 0.0461296f
c3 4 VSS 0.00471071f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1207 $X2=0.1890 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1150 $X2=0.1890 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1150 $X2=0.1890 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AOI332xp33_ASAP7_75t_R%C2 VSS 6 3 4 1
c1 1 VSS 0.00794248f
c2 3 VSS 0.0466528f
c3 4 VSS 0.00501592f
r1 7 8 3.43955 $w=1.3e-08 $l=1.48e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1202 $X2=0.4050 $Y2=0.1350
r2 6 7 1.45744 $w=1.3e-08 $l=6.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1140 $X2=0.4050 $Y2=0.1202
r3 6 4 5.18847 $w=1.3e-08 $l=2.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1140 $X2=0.4050 $Y2=0.0917
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
.ends

.subckt PM_AOI332xp33_ASAP7_75t_R%B1 VSS 6 3 1 4
c1 1 VSS 0.00831977f
c2 3 VSS 0.00945592f
c3 4 VSS 0.00522092f
r1 7 8 3.20636 $w=1.3e-08 $l=1.38e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1212 $X2=0.2430 $Y2=0.1350
r2 6 7 1.22425 $w=1.3e-08 $l=5.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1160 $X2=0.2430 $Y2=0.1212
r3 6 4 5.42166 $w=1.3e-08 $l=2.33e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1160 $X2=0.2430 $Y2=0.0927
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AOI332xp33_ASAP7_75t_R%B3 VSS 6 3 1 4
c1 1 VSS 0.00796311f
c2 3 VSS 0.0468132f
c3 4 VSS 0.00514742f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1207 $X2=0.3510 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1150 $X2=0.3510 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1150 $X2=0.3510 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
.ends

.subckt PM_AOI332xp33_ASAP7_75t_R%Y VSS 39 20 21 43 51 52 13 10 1 14 2 12 3 15
+ 11 17
c1 1 VSS 0.00660589f
c2 2 VSS 0.00277208f
c3 3 VSS 0.00550687f
c4 10 VSS 0.00341067f
c5 11 VSS 0.00269163f
c6 12 VSS 0.00215412f
c7 13 VSS 0.0288986f
c8 14 VSS 0.000743886f
c9 15 VSS 0.00209502f
c10 16 VSS 0.00275231f
c11 17 VSS 0.000781121f
r1 52 50 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r2 2 50 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r3 12 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r4 51 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r5 2 47 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.1980
r6 47 48 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.1980 $X2=0.4455 $Y2=0.1980
r7 45 48 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1980 $X2=0.4455 $Y2=0.1980
r8 44 45 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.4850
+ $Y=0.1980 $X2=0.4590 $Y2=0.1980
r9 14 17 0.682785 $w=1.75e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5030
+ $Y=0.1980 $X2=0.5130 $Y2=0.1980
r10 14 44 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5030
+ $Y=0.1980 $X2=0.4850 $Y2=0.1980
r11 17 41 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1980 $X2=0.5130 $Y2=0.1765
r12 11 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0675 $X2=0.4840 $Y2=0.0675
r13 43 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4715 $Y2=0.0675
r14 40 41 7.17059 $w=1.3e-08 $l=3.08e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1457 $X2=0.5130 $Y2=0.1765
r15 39 40 4.37231 $w=1.3e-08 $l=1.87e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1270 $X2=0.5130 $Y2=0.1457
r16 39 38 6.70421 $w=1.3e-08 $l=2.88e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1270 $X2=0.5130 $Y2=0.0982
r17 15 16 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.0575 $X2=0.5130 $Y2=0.0360
r18 15 38 9.50248 $w=1.3e-08 $l=4.07e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0575 $X2=0.5130 $Y2=0.0982
r19 3 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0675
+ $X2=0.4860 $Y2=0.0360
r20 16 37 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.0360 $X2=0.4995 $Y2=0.0360
r21 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.0360 $X2=0.4995 $Y2=0.0360
r22 35 36 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4725
+ $Y=0.0360 $X2=0.4860 $Y2=0.0360
r23 34 35 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0360 $X2=0.4725 $Y2=0.0360
r24 33 34 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.4335
+ $Y=0.0360 $X2=0.4590 $Y2=0.0360
r25 32 33 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4155
+ $Y=0.0360 $X2=0.4335 $Y2=0.0360
r26 31 32 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0360 $X2=0.4155 $Y2=0.0360
r27 30 31 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0360 $X2=0.4050 $Y2=0.0360
r28 29 30 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r29 28 29 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.3405
+ $Y=0.0360 $X2=0.3510 $Y2=0.0360
r30 27 28 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3225
+ $Y=0.0360 $X2=0.3405 $Y2=0.0360
r31 26 27 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.3225 $Y2=0.0360
r32 25 26 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.2970 $Y2=0.0360
r33 24 25 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r34 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r35 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.2295 $Y2=0.0360
r36 13 22 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2040
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r37 1 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0675
+ $X2=0.2160 $Y2=0.0360
r38 21 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r39 1 19 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r40 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r41 20 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2015 $Y2=0.0675
.ends

.subckt PM_AOI332xp33_ASAP7_75t_R%NET030 VSS 16 17 32 33 35 10 1 11 2 12 3 13
c1 1 VSS 0.00474593f
c2 2 VSS 0.00413884f
c3 3 VSS 0.00522703f
c4 10 VSS 0.00222326f
c5 11 VSS 0.00220175f
c6 12 VSS 0.00228512f
c7 13 VSS 0.0205709f
r1 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4840 $Y2=0.2025
r2 35 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r3 33 31 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r4 2 31 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r5 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3780 $Y2=0.2025
r6 32 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r7 3 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2025
+ $X2=0.4860 $Y2=0.2340
r8 2 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.2340
r9 27 28 9.0944 $w=1.3e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4470
+ $Y=0.2340 $X2=0.4860 $Y2=0.2340
r10 26 27 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4155
+ $Y=0.2340 $X2=0.4470 $Y2=0.2340
r11 25 26 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.2340 $X2=0.4155 $Y2=0.2340
r12 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3915
+ $Y=0.2340 $X2=0.4050 $Y2=0.2340
r13 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r14 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3645
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r15 21 22 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.2340 $X2=0.3645 $Y2=0.2340
r16 20 21 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.3405
+ $Y=0.2340 $X2=0.3510 $Y2=0.2340
r17 19 20 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3090
+ $Y=0.2340 $X2=0.3405 $Y2=0.2340
r18 18 19 9.0944 $w=1.3e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.3090 $Y2=0.2340
r19 13 18 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2575
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r20 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.2340
r21 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r22 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r23 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r24 16 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
.ends


*
.SUBCKT AOI332xp33_ASAP7_75t_R VSS VDD A3 A2 A1 B1 B2 B3 C2 C1 Y
*
* VSS VSS
* VDD VDD
* A3 A3
* A2 A2
* A1 A1
* B1 B1
* B2 B2
* B3 B3
* C2 C2
* C1 C1
* Y Y
*
*

MM3 N_MM3_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM14 N_MM14_d N_MM9_g N_MM14_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM12 N_MM12_d N_MM6_g N_MM12_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 N_MM11_d N_MM5_g N_MM11_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM16 N_MM16_d N_MM0_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM17 N_MM17_d N_MM1_g N_MM17_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM6_g N_MM6_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g N_MM4_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM0_g N_MM0_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AOI332xp33_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AOI332xp33_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AOI332xp33_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_AOI332xp33_ASAP7_75t_R%noxref_20
cc_1 N_noxref_20_1 N_MM3_g 0.0016098f
cc_2 N_noxref_20_1 N_noxref_19_1 0.00179267f
x_PM_AOI332xp33_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_AOI332xp33_ASAP7_75t_R%noxref_19
cc_3 N_noxref_19_1 N_MM3_g 0.00165616f
x_PM_AOI332xp33_ASAP7_75t_R%NET061 VSS N_MM16_d N_MM17_s N_NET061_1
+ PM_AOI332xp33_ASAP7_75t_R%NET061
cc_4 N_NET061_1 N_MM0_g 0.0172826f
cc_5 N_NET061_1 N_MM1_g 0.0171848f
x_PM_AOI332xp33_ASAP7_75t_R%NET064 VSS N_MM11_s N_MM10_d N_NET064_1
+ PM_AOI332xp33_ASAP7_75t_R%NET064
cc_6 N_NET064_1 N_MM5_g 0.0173954f
cc_7 N_NET064_1 N_MM4_g 0.0173009f
x_PM_AOI332xp33_ASAP7_75t_R%NET063 VSS N_MM12_s N_MM11_d N_NET063_1
+ PM_AOI332xp33_ASAP7_75t_R%NET063
cc_8 N_NET063_1 N_MM6_g 0.0173774f
cc_9 N_NET063_1 N_MM5_g 0.0173005f
x_PM_AOI332xp33_ASAP7_75t_R%NET25 VSS N_MM3_d N_MM2_s N_NET25_1
+ PM_AOI332xp33_ASAP7_75t_R%NET25
cc_10 N_NET25_1 N_MM3_g 0.0173493f
cc_11 N_NET25_1 N_MM2_g 0.0173018f
x_PM_AOI332xp33_ASAP7_75t_R%NET26 VSS N_MM2_d N_MM14_s N_NET26_1
+ PM_AOI332xp33_ASAP7_75t_R%NET26
cc_12 N_NET26_1 N_MM2_g 0.0172993f
cc_13 N_NET26_1 N_MM9_g 0.0171696f
x_PM_AOI332xp33_ASAP7_75t_R%A2 VSS A2 N_MM2_g N_A2_1 N_A2_4
+ PM_AOI332xp33_ASAP7_75t_R%A2
cc_14 N_A2_1 N_A3_1 0.00131187f
cc_15 N_A2_4 N_A3_4 0.00522118f
cc_16 N_MM2_g N_MM3_g 0.00631375f
x_PM_AOI332xp33_ASAP7_75t_R%A3 VSS A3 N_MM3_g N_A3_1 N_A3_4
+ PM_AOI332xp33_ASAP7_75t_R%A3
x_PM_AOI332xp33_ASAP7_75t_R%NET031 VSS N_MM9_d N_MM6_s N_MM7_d N_MM8_d N_MM5_s
+ N_MM4_s N_NET031_13 N_NET031_1 N_NET031_10 N_NET031_2 N_NET031_11 N_NET031_12
+ N_NET031_3 PM_AOI332xp33_ASAP7_75t_R%NET031
cc_17 N_NET031_13 N_A3_4 0.000740175f
cc_18 N_NET031_1 N_MM3_g 0.000905885f
cc_19 N_NET031_1 N_A3_4 0.000932741f
cc_20 N_NET031_10 N_MM3_g 0.0341497f
cc_21 N_NET031_10 N_A2_1 0.000728683f
cc_22 N_NET031_1 N_MM2_g 0.000878219f
cc_23 N_NET031_13 N_A2_4 0.00124067f
cc_24 N_NET031_1 N_A2_4 0.0012531f
cc_25 N_NET031_10 N_MM2_g 0.033517f
cc_26 N_NET031_2 N_MM9_g 0.000868745f
cc_27 N_NET031_2 N_A1_4 0.00126358f
cc_28 N_NET031_13 N_A1_4 0.001272f
cc_29 N_NET031_11 N_MM9_g 0.0342411f
cc_30 N_NET031_11 N_B1_1 0.000859761f
cc_31 N_NET031_2 N_MM6_g 0.000866671f
cc_32 N_NET031_13 N_B1_4 0.00125732f
cc_33 N_NET031_2 N_B1_4 0.00127528f
cc_34 N_NET031_11 N_MM6_g 0.0333845f
cc_35 N_NET031_12 N_B2_1 0.00076933f
cc_36 N_NET031_3 N_MM5_g 0.000868692f
cc_37 N_NET031_13 N_B2_4 0.00120989f
cc_38 N_NET031_3 N_B2_4 0.00121f
cc_39 N_NET031_12 N_MM5_g 0.0335112f
cc_40 N_NET031_12 N_B3_1 0.000745538f
cc_41 N_NET031_3 N_B3_4 0.000761135f
cc_42 N_NET031_3 N_MM4_g 0.0008915f
cc_43 N_NET031_12 N_MM4_g 0.033865f
x_PM_AOI332xp33_ASAP7_75t_R%B2 VSS B2 N_MM5_g N_B2_1 N_B2_4
+ PM_AOI332xp33_ASAP7_75t_R%B2
cc_44 N_B2_1 N_B1_1 0.00137943f
cc_45 N_B2_4 N_B1_4 0.00331567f
cc_46 N_MM5_g N_MM6_g 0.00607119f
x_PM_AOI332xp33_ASAP7_75t_R%C1 VSS C1 N_MM1_g N_C1_1 N_C1_4
+ PM_AOI332xp33_ASAP7_75t_R%C1
cc_47 N_C1_1 N_C2_1 0.00128998f
cc_48 N_C1_4 N_C2_4 0.0033851f
cc_49 N_MM1_g N_MM0_g 0.00587839f
x_PM_AOI332xp33_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_AOI332xp33_ASAP7_75t_R%noxref_21
cc_50 N_noxref_21_1 N_MM1_g 0.00145974f
cc_51 N_noxref_21_1 N_NET030_12 0.000472023f
cc_52 N_noxref_21_1 N_Y_11 0.0372307f
x_PM_AOI332xp33_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_AOI332xp33_ASAP7_75t_R%noxref_22
cc_53 N_noxref_22_1 N_MM1_g 0.0014506f
cc_54 N_noxref_22_1 N_NET030_12 0.035976f
cc_55 N_noxref_22_1 N_Y_12 0.00120302f
cc_56 N_noxref_22_1 N_noxref_21_1 0.00176539f
x_PM_AOI332xp33_ASAP7_75t_R%A1 VSS A1 N_MM9_g N_A1_1 N_A1_4
+ PM_AOI332xp33_ASAP7_75t_R%A1
cc_57 N_A1_1 N_A2_1 0.00129658f
cc_58 N_A1_4 N_A2_4 0.00399157f
cc_59 N_MM9_g N_MM2_g 0.0061957f
x_PM_AOI332xp33_ASAP7_75t_R%C2 VSS C2 N_MM0_g N_C2_4 N_C2_1
+ PM_AOI332xp33_ASAP7_75t_R%C2
cc_60 N_C2_4 N_B3_1 0.000936951f
cc_61 N_MM0_g N_MM4_g 0.00326796f
cc_62 N_C2_4 N_B3_4 0.00413537f
x_PM_AOI332xp33_ASAP7_75t_R%B1 VSS B1 N_MM6_g N_B1_1 N_B1_4
+ PM_AOI332xp33_ASAP7_75t_R%B1
cc_63 N_B1_1 N_MM9_g 0.000920505f
cc_64 N_B1_4 N_A1_4 0.00319167f
cc_65 N_MM6_g N_MM9_g 0.00400514f
x_PM_AOI332xp33_ASAP7_75t_R%B3 VSS B3 N_MM4_g N_B3_1 N_B3_4
+ PM_AOI332xp33_ASAP7_75t_R%B3
cc_66 N_B3_1 N_B2_1 0.00127319f
cc_67 N_B3_4 N_B2_4 0.0033943f
cc_68 N_MM4_g N_MM5_g 0.0059838f
x_PM_AOI332xp33_ASAP7_75t_R%Y VSS Y N_MM14_d N_MM12_d N_MM17_d N_MM0_d N_MM1_d
+ N_Y_13 N_Y_10 N_Y_1 N_Y_14 N_Y_2 N_Y_12 N_Y_3 N_Y_15 N_Y_11 N_Y_17
+ PM_AOI332xp33_ASAP7_75t_R%Y
cc_69 N_Y_13 N_MM9_g 0.000555887f
cc_70 N_Y_10 N_A1_1 0.000743479f
cc_71 N_Y_1 N_A1_4 0.00120663f
cc_72 N_Y_1 N_MM9_g 0.00155586f
cc_73 N_Y_10 N_MM9_g 0.0350735f
cc_74 N_Y_10 N_B1_1 0.000884148f
cc_75 N_Y_13 N_B1_4 0.00119597f
cc_76 N_Y_1 N_MM6_g 0.00153658f
cc_77 N_Y_1 N_B1_4 0.00169128f
cc_78 N_Y_10 N_MM6_g 0.0349863f
cc_79 N_Y_13 N_B2_4 0.00374334f
cc_80 N_Y_13 N_B3_4 0.00317069f
cc_81 N_Y_14 N_C2_4 0.000573905f
cc_82 N_Y_2 N_MM0_g 0.000924715f
cc_83 N_Y_12 N_C2_1 0.000937815f
cc_84 N_Y_13 N_C2_4 0.00129287f
cc_85 N_Y_2 N_C2_4 0.00213673f
cc_86 N_Y_12 N_MM0_g 0.0353595f
cc_87 N_Y_2 N_C1_1 0.000897217f
cc_88 N_Y_2 N_MM1_g 0.000910889f
cc_89 N_Y_14 N_C1_4 0.00102064f
cc_90 N_Y_13 N_C1_4 0.00115977f
cc_91 N_Y_3 N_MM1_g 0.00165258f
cc_92 N_Y_12 N_C1_1 0.001697f
cc_93 N_Y_12 N_MM1_g 0.0149906f
cc_94 N_Y_15 N_C1_4 0.00656763f
cc_95 N_Y_11 N_MM1_g 0.054248f
cc_96 N_Y_12 N_NET030_11 0.00168256f
cc_97 N_Y_15 N_NET030_3 0.000718086f
cc_98 N_Y_17 N_NET030_13 0.000730726f
cc_99 N_Y_12 N_NET030_12 0.000767056f
cc_100 N_Y_2 N_NET030_13 0.000792851f
cc_101 N_Y_2 N_NET030_3 0.00253167f
cc_102 N_Y_2 N_NET030_2 0.00416219f
cc_103 N_Y_14 N_NET030_13 0.00966408f
x_PM_AOI332xp33_ASAP7_75t_R%NET030 VSS N_MM6_d N_MM5_d N_MM4_d N_MM0_s N_MM1_s
+ N_NET030_10 N_NET030_1 N_NET030_11 N_NET030_2 N_NET030_12 N_NET030_3
+ N_NET030_13 PM_AOI332xp33_ASAP7_75t_R%NET030
cc_104 N_NET030_10 N_B1_1 0.000787892f
cc_105 N_NET030_1 N_MM6_g 0.000913491f
cc_106 N_NET030_10 N_MM6_g 0.0338702f
cc_107 N_NET030_10 N_B2_1 0.000763427f
cc_108 N_NET030_1 N_MM5_g 0.000912616f
cc_109 N_NET030_10 N_MM5_g 0.0340058f
cc_110 N_NET030_11 N_B3_1 0.000728962f
cc_111 N_NET030_2 N_MM4_g 0.000970045f
cc_112 N_NET030_11 N_MM4_g 0.0343915f
cc_113 N_NET030_11 N_C2_1 0.000810352f
cc_114 N_NET030_2 N_MM0_g 0.000948144f
cc_115 N_NET030_11 N_MM0_g 0.0343374f
cc_116 N_NET030_12 N_C1_1 0.000739059f
cc_117 N_NET030_3 N_MM1_g 0.00101479f
cc_118 N_NET030_12 N_MM1_g 0.0342352f
cc_119 N_NET030_10 N_NET031_13 0.000553082f
cc_120 N_NET030_1 N_NET031_13 0.00068195f
cc_121 N_NET030_13 N_NET031_3 0.000748148f
cc_122 N_NET030_10 N_NET031_12 0.00111317f
cc_123 N_NET030_10 N_NET031_11 0.00111785f
cc_124 N_NET030_2 N_NET031_3 0.00133187f
cc_125 N_NET030_1 N_NET031_3 0.00275017f
cc_126 N_NET030_1 N_NET031_2 0.00423689f
cc_127 N_NET030_13 N_NET031_13 0.0100749f
*END of AOI332xp33_ASAP7_75t_R.pxi
.ENDS
** Design:	AOI333xp33_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AOI333xp33_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AOI333xp33_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AOI333xp33_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.0429131f
.ends

.subckt PM_AOI333xp33_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.0429204f
.ends

.subckt PM_AOI333xp33_ASAP7_75t_R%NET25 VSS 2 3 1
c1 1 VSS 0.00097564f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4320 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4320 $Y2=0.0675
.ends

.subckt PM_AOI333xp33_ASAP7_75t_R%NET063 VSS 2 3 1
c1 1 VSS 0.0010075f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2700 $Y2=0.0675
.ends

.subckt PM_AOI333xp33_ASAP7_75t_R%NET064 VSS 2 3 1
c1 1 VSS 0.000994435f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3240 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3240 $Y2=0.0675
.ends

.subckt PM_AOI333xp33_ASAP7_75t_R%NET062 VSS 2 3 1
c1 1 VSS 0.00094816f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_AOI333xp33_ASAP7_75t_R%NET061 VSS 2 3 1
c1 1 VSS 0.0009491f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_AOI333xp33_ASAP7_75t_R%NET26 VSS 2 3 1
c1 1 VSS 0.000963161f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4860 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0675 $X2=0.4860 $Y2=0.0675
.ends

.subckt PM_AOI333xp33_ASAP7_75t_R%C2 VSS 6 3 1 4
c1 1 VSS 0.00706885f
c2 3 VSS 0.047383f
c3 4 VSS 0.00831352f
r1 7 8 3.20636 $w=1.3e-08 $l=1.38e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1212 $X2=0.1350 $Y2=0.1350
r2 6 7 1.22425 $w=1.3e-08 $l=5.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1160 $X2=0.1350 $Y2=0.1212
r3 6 4 5.42166 $w=1.3e-08 $l=2.33e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1160 $X2=0.1350 $Y2=0.0927
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AOI333xp33_ASAP7_75t_R%C3 VSS 6 3 1 4
c1 1 VSS 0.00556171f
c2 3 VSS 0.0820909f
c3 4 VSS 0.0162915f
r1 7 8 3.43955 $w=1.3e-08 $l=1.48e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1202 $X2=0.0810 $Y2=0.1350
r2 6 7 1.45744 $w=1.3e-08 $l=6.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1140 $X2=0.0810 $Y2=0.1202
r3 6 4 9.38589 $w=1.3e-08 $l=4.03e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1140 $X2=0.0810 $Y2=0.0737
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AOI333xp33_ASAP7_75t_R%NET031 VSS 16 17 36 37 40 41 13 1 10 2 11 12 3
c1 1 VSS 0.00890016f
c2 2 VSS 0.00592489f
c3 3 VSS 0.002939f
c4 10 VSS 0.00453025f
c5 11 VSS 0.00334498f
c6 12 VSS 0.00214177f
c7 13 VSS 0.00798523f
r1 41 39 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r2 3 39 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r3 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r4 40 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r5 37 35 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r6 2 35 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r7 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r8 36 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r9 3 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.1980
r10 2 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.1980
r11 31 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3105
+ $Y=0.1980 $X2=0.3240 $Y2=0.1980
r12 30 31 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1980 $X2=0.3105 $Y2=0.1980
r13 29 30 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2710
+ $Y=0.1980 $X2=0.2970 $Y2=0.1980
r14 28 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2530
+ $Y=0.1980 $X2=0.2710 $Y2=0.1980
r15 27 28 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1980 $X2=0.2530 $Y2=0.1980
r16 26 27 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.1980 $X2=0.2430 $Y2=0.1980
r17 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1980 $X2=0.2295 $Y2=0.1980
r18 24 25 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2040
+ $Y=0.1980 $X2=0.2160 $Y2=0.1980
r19 23 24 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1995
+ $Y=0.1980 $X2=0.2040 $Y2=0.1980
r20 22 23 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1980 $X2=0.1995 $Y2=0.1980
r21 21 22 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.1980 $X2=0.1890 $Y2=0.1980
r22 20 21 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1980 $X2=0.1620 $Y2=0.1980
r23 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1215
+ $Y=0.1980 $X2=0.1350 $Y2=0.1980
r24 18 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.1980 $X2=0.1215 $Y2=0.1980
r25 13 18 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0965
+ $Y=0.1980 $X2=0.1080 $Y2=0.1980
r26 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.1980
r27 16 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r28 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r29 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r30 17 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
.ends

.subckt PM_AOI333xp33_ASAP7_75t_R%B1 VSS 6 3 1 4
c1 1 VSS 0.00799123f
c2 3 VSS 0.00927167f
c3 4 VSS 0.00507981f
r1 7 8 3.20636 $w=1.3e-08 $l=1.38e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1212 $X2=0.2430 $Y2=0.1350
r2 6 7 1.22425 $w=1.3e-08 $l=5.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1160 $X2=0.2430 $Y2=0.1212
r3 6 4 5.42166 $w=1.3e-08 $l=2.33e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1160 $X2=0.2430 $Y2=0.0927
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AOI333xp33_ASAP7_75t_R%B2 VSS 6 3 1 4
c1 1 VSS 0.00727745f
c2 3 VSS 0.00976631f
c3 4 VSS 0.00483378f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1207 $X2=0.2970 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1150 $X2=0.2970 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1150 $X2=0.2970 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_AOI333xp33_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.00530964f
.ends

.subckt PM_AOI333xp33_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.00525007f
.ends

.subckt PM_AOI333xp33_ASAP7_75t_R%C1 VSS 6 3 1 4
c1 1 VSS 0.00769914f
c2 3 VSS 0.0460391f
c3 4 VSS 0.00463495f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1207 $X2=0.1890 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1150 $X2=0.1890 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1150 $X2=0.1890 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AOI333xp33_ASAP7_75t_R%A3 VSS 6 3 4 1
c1 1 VSS 0.00781188f
c2 3 VSS 0.0466568f
c3 4 VSS 0.00511136f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1207 $X2=0.4050 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1150 $X2=0.4050 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1150 $X2=0.4050 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
.ends

.subckt PM_AOI333xp33_ASAP7_75t_R%A1 VSS 6 3 1 4
c1 1 VSS 0.00750923f
c2 3 VSS 0.00878381f
c3 4 VSS 0.00450337f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1207 $X2=0.5130 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1150 $X2=0.5130 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1150 $X2=0.5130 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.1350
+ $X2=0.5130 $Y2=0.1350
.ends

.subckt PM_AOI333xp33_ASAP7_75t_R%B3 VSS 6 3 1 4
c1 1 VSS 0.0082162f
c2 3 VSS 0.0468067f
c3 4 VSS 0.00511523f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1207 $X2=0.3510 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1150 $X2=0.3510 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1150 $X2=0.3510 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
.ends

.subckt PM_AOI333xp33_ASAP7_75t_R%A2 VSS 6 3 1 4
c1 1 VSS 0.00654509f
c2 3 VSS 0.00943883f
c3 4 VSS 0.00427603f
r1 7 8 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1207 $X2=0.4590 $Y2=0.1350
r2 6 7 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1150 $X2=0.4590 $Y2=0.1207
r3 6 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1150 $X2=0.4590 $Y2=0.0922
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1350
+ $X2=0.4590 $Y2=0.1350
.ends

.subckt PM_AOI333xp33_ASAP7_75t_R%Y VSS 44 24 25 48 60 63 64 17 13 1 18 2 15 16
+ 4 3 19 14
c1 1 VSS 0.00665828f
c2 2 VSS 0.00292914f
c3 3 VSS 0.00548721f
c4 4 VSS 0.00406235f
c5 13 VSS 0.00345366f
c6 14 VSS 0.00268912f
c7 15 VSS 0.00220158f
c8 16 VSS 0.00235393f
c9 17 VSS 0.0349896f
c10 18 VSS 0.00177758f
c11 19 VSS 0.00226604f
c12 20 VSS 0.00288086f
c13 21 VSS 0.00112078f
r1 64 62 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r2 2 62 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r3 15 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r4 63 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r5 16 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.2025 $X2=0.5380 $Y2=0.2025
r6 60 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.2025 $X2=0.5255 $Y2=0.2025
r7 2 56 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.1980
r8 4 49 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.2025
+ $X2=0.5400 $Y2=0.1980
r9 56 57 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.1980 $X2=0.4455 $Y2=0.1980
r10 54 57 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1980 $X2=0.4455 $Y2=0.1980
r11 53 54 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.1980 $X2=0.4590 $Y2=0.1980
r12 52 53 5.47996 $w=1.3e-08 $l=2.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5095
+ $Y=0.1980 $X2=0.4860 $Y2=0.1980
r13 51 52 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5185
+ $Y=0.1980 $X2=0.5095 $Y2=0.1980
r14 49 50 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1980 $X2=0.5535 $Y2=0.1980
r15 18 49 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5265
+ $Y=0.1980 $X2=0.5400 $Y2=0.1980
r16 18 51 1.86552 $w=1.3e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.5265
+ $Y=0.1980 $X2=0.5185 $Y2=0.1980
r17 21 46 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.1980 $X2=0.5670 $Y2=0.1765
r18 21 50 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.1980 $X2=0.5535 $Y2=0.1980
r19 14 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.0675 $X2=0.5380 $Y2=0.0675
r20 48 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.0675 $X2=0.5255 $Y2=0.0675
r21 45 46 7.17059 $w=1.3e-08 $l=3.08e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1457 $X2=0.5670 $Y2=0.1765
r22 44 45 4.37231 $w=1.3e-08 $l=1.87e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1270 $X2=0.5670 $Y2=0.1457
r23 44 43 6.70421 $w=1.3e-08 $l=2.88e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1270 $X2=0.5670 $Y2=0.0982
r24 19 20 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.0575 $X2=0.5670 $Y2=0.0360
r25 19 43 9.50248 $w=1.3e-08 $l=4.07e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0575 $X2=0.5670 $Y2=0.0982
r26 3 41 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.0675
+ $X2=0.5400 $Y2=0.0360
r27 20 42 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.0360 $X2=0.5535 $Y2=0.0360
r28 41 42 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.0360 $X2=0.5535 $Y2=0.0360
r29 40 41 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5265
+ $Y=0.0360 $X2=0.5400 $Y2=0.0360
r30 39 40 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0360 $X2=0.5265 $Y2=0.0360
r31 38 39 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.0360 $X2=0.5130 $Y2=0.0360
r32 37 38 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0360 $X2=0.4860 $Y2=0.0360
r33 36 37 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4590 $Y2=0.0360
r34 35 36 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r35 34 35 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0360 $X2=0.4050 $Y2=0.0360
r36 33 34 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r37 32 33 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3410
+ $Y=0.0360 $X2=0.3510 $Y2=0.0360
r38 31 32 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3230
+ $Y=0.0360 $X2=0.3410 $Y2=0.0360
r39 30 31 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.3230 $Y2=0.0360
r40 29 30 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.2970 $Y2=0.0360
r41 28 29 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r42 27 28 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r43 26 27 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.2295 $Y2=0.0360
r44 17 26 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2040
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r45 1 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0675
+ $X2=0.2160 $Y2=0.0360
r46 25 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r47 1 23 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r48 13 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r49 24 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2015 $Y2=0.0675
.ends

.subckt PM_AOI333xp33_ASAP7_75t_R%NET030 VSS 16 17 31 32 35 36 1 10 11 2 12 3 13
c1 1 VSS 0.0046369f
c2 2 VSS 0.00427318f
c3 3 VSS 0.00444962f
c4 10 VSS 0.00214609f
c5 11 VSS 0.00213438f
c6 12 VSS 0.00214736f
c7 13 VSS 0.0217463f
r1 36 34 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r2 3 34 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r3 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4860 $Y2=0.2025
r4 35 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r5 32 30 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r6 2 30 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r7 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3780 $Y2=0.2025
r8 31 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r9 3 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2025
+ $X2=0.4860 $Y2=0.2340
r10 2 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.2340
r11 26 27 9.56078 $w=1.3e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4450
+ $Y=0.2340 $X2=0.4860 $Y2=0.2340
r12 25 26 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4045
+ $Y=0.2340 $X2=0.4450 $Y2=0.2340
r13 24 25 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.3915
+ $Y=0.2340 $X2=0.4045 $Y2=0.2340
r14 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r15 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3645
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r16 21 22 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.2340 $X2=0.3645 $Y2=0.2340
r17 20 21 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3410
+ $Y=0.2340 $X2=0.3510 $Y2=0.2340
r18 19 20 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3095
+ $Y=0.2340 $X2=0.3410 $Y2=0.2340
r19 18 19 9.211 $w=1.3e-08 $l=3.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.3095 $Y2=0.2340
r20 13 18 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2575
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r21 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.2340
r22 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r23 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r24 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r25 16 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
.ends


*
.SUBCKT AOI333xp33_ASAP7_75t_R VSS VDD C3 C2 C1 B1 B2 B3 A3 A2 A1 Y
*
* VSS VSS
* VDD VDD
* C3 C3
* C2 C2
* C1 C1
* B1 B1
* B2 B2
* B3 B3
* A3 A3
* A2 A2
* A1 A1
* Y Y
*
*

MM13 N_MM13_d N_MM13_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM16 N_MM16_d N_MM8_g N_MM16_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM17 N_MM17_d N_MM9_g N_MM17_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM12 N_MM12_d N_MM6_g N_MM12_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 N_MM11_d N_MM5_g N_MM11_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM15_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM0_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM14 N_MM14_d N_MM1_g N_MM14_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM13_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM8_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM6_g N_MM6_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g N_MM4_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM15 N_MM15_d N_MM15_g N_MM15_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM0_g N_MM0_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AOI333xp33_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AOI333xp33_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AOI333xp33_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_AOI333xp33_ASAP7_75t_R%noxref_21
cc_1 N_noxref_21_1 N_MM13_g 0.00165685f
x_PM_AOI333xp33_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_AOI333xp33_ASAP7_75t_R%noxref_22
cc_2 N_noxref_22_1 N_MM13_g 0.00161594f
cc_3 N_noxref_22_1 N_noxref_21_1 0.00179488f
x_PM_AOI333xp33_ASAP7_75t_R%NET25 VSS N_MM3_d N_MM2_s N_NET25_1
+ PM_AOI333xp33_ASAP7_75t_R%NET25
cc_4 N_NET25_1 N_MM15_g 0.017357f
cc_5 N_NET25_1 N_MM0_g 0.0173559f
x_PM_AOI333xp33_ASAP7_75t_R%NET063 VSS N_MM12_s N_MM11_d N_NET063_1
+ PM_AOI333xp33_ASAP7_75t_R%NET063
cc_6 N_NET063_1 N_MM6_g 0.0173808f
cc_7 N_NET063_1 N_MM5_g 0.0173002f
x_PM_AOI333xp33_ASAP7_75t_R%NET064 VSS N_MM11_s N_MM10_d N_NET064_1
+ PM_AOI333xp33_ASAP7_75t_R%NET064
cc_8 N_NET064_1 N_MM5_g 0.0173898f
cc_9 N_NET064_1 N_MM4_g 0.0173037f
x_PM_AOI333xp33_ASAP7_75t_R%NET062 VSS N_MM13_d N_MM16_s N_NET062_1
+ PM_AOI333xp33_ASAP7_75t_R%NET062
cc_10 N_NET062_1 N_MM13_g 0.0173528f
cc_11 N_NET062_1 N_MM8_g 0.0172973f
x_PM_AOI333xp33_ASAP7_75t_R%NET061 VSS N_MM16_d N_MM17_s N_NET061_1
+ PM_AOI333xp33_ASAP7_75t_R%NET061
cc_12 N_NET061_1 N_MM8_g 0.0172958f
cc_13 N_NET061_1 N_MM9_g 0.0171727f
x_PM_AOI333xp33_ASAP7_75t_R%NET26 VSS N_MM2_d N_MM14_s N_NET26_1
+ PM_AOI333xp33_ASAP7_75t_R%NET26
cc_14 N_NET26_1 N_MM0_g 0.0173432f
cc_15 N_NET26_1 N_MM1_g 0.0171735f
x_PM_AOI333xp33_ASAP7_75t_R%C2 VSS C2 N_MM8_g N_C2_1 N_C2_4
+ PM_AOI333xp33_ASAP7_75t_R%C2
cc_16 N_C2_1 N_C3_1 0.00131196f
cc_17 N_C2_4 N_C3_4 0.00509506f
cc_18 N_MM8_g N_MM13_g 0.0063069f
x_PM_AOI333xp33_ASAP7_75t_R%C3 VSS C3 N_MM13_g N_C3_1 N_C3_4
+ PM_AOI333xp33_ASAP7_75t_R%C3
x_PM_AOI333xp33_ASAP7_75t_R%NET031 VSS N_MM8_d N_MM7_d N_MM9_d N_MM6_s N_MM5_s
+ N_MM4_s N_NET031_13 N_NET031_1 N_NET031_10 N_NET031_2 N_NET031_11 N_NET031_12
+ N_NET031_3 PM_AOI333xp33_ASAP7_75t_R%NET031
cc_19 N_NET031_13 N_C3_4 0.000720128f
cc_20 N_NET031_1 N_C3_4 0.000886389f
cc_21 N_NET031_1 N_MM13_g 0.000908098f
cc_22 N_NET031_10 N_MM13_g 0.0342351f
cc_23 N_NET031_10 N_C2_1 0.000730203f
cc_24 N_NET031_1 N_MM8_g 0.000879804f
cc_25 N_NET031_13 N_C2_4 0.00127179f
cc_26 N_NET031_1 N_C2_4 0.00127487f
cc_27 N_NET031_10 N_MM8_g 0.0336015f
cc_28 N_NET031_2 N_MM9_g 0.000870758f
cc_29 N_NET031_2 N_C1_4 0.00127784f
cc_30 N_NET031_13 N_C1_4 0.00128142f
cc_31 N_NET031_11 N_MM9_g 0.0343202f
cc_32 N_NET031_11 N_B1_1 0.00060053f
cc_33 N_NET031_2 N_MM6_g 0.000868679f
cc_34 N_NET031_13 N_B1_4 0.0012625f
cc_35 N_NET031_2 N_B1_4 0.00127847f
cc_36 N_NET031_11 N_MM6_g 0.0334625f
cc_37 N_NET031_12 N_B2_1 0.000755632f
cc_38 N_NET031_3 N_MM5_g 0.000882701f
cc_39 N_NET031_3 N_B2_4 0.00119617f
cc_40 N_NET031_13 N_B2_4 0.00122195f
cc_41 N_NET031_12 N_MM5_g 0.0335829f
cc_42 N_NET031_13 N_B3_4 0.000642298f
cc_43 N_NET031_3 N_B3_4 0.000804455f
cc_44 N_NET031_3 N_MM4_g 0.000899068f
cc_45 N_NET031_12 N_MM4_g 0.0339006f
x_PM_AOI333xp33_ASAP7_75t_R%B1 VSS B1 N_MM6_g N_B1_1 N_B1_4
+ PM_AOI333xp33_ASAP7_75t_R%B1
cc_46 N_B1_1 N_MM9_g 0.000863321f
cc_47 N_B1_4 N_C1_4 0.00319363f
cc_48 N_MM6_g N_MM9_g 0.0040053f
x_PM_AOI333xp33_ASAP7_75t_R%B2 VSS B2 N_MM5_g N_B2_1 N_B2_4
+ PM_AOI333xp33_ASAP7_75t_R%B2
cc_49 N_B2_1 N_B1_1 0.00127625f
cc_50 N_B2_4 N_B1_4 0.00332606f
cc_51 N_MM5_g N_MM6_g 0.00607082f
x_PM_AOI333xp33_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_AOI333xp33_ASAP7_75t_R%noxref_23
cc_52 N_noxref_23_1 N_MM1_g 0.00145691f
cc_53 N_noxref_23_1 N_Y_3 0.000501472f
cc_54 N_noxref_23_1 N_Y_14 0.0374468f
x_PM_AOI333xp33_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_AOI333xp33_ASAP7_75t_R%noxref_24
cc_55 N_noxref_24_1 N_MM1_g 0.00144606f
cc_56 N_noxref_24_1 N_Y_4 0.00049902f
cc_57 N_noxref_24_1 N_Y_16 0.0375002f
cc_58 N_noxref_24_1 N_noxref_23_1 0.00177342f
x_PM_AOI333xp33_ASAP7_75t_R%C1 VSS C1 N_MM9_g N_C1_1 N_C1_4
+ PM_AOI333xp33_ASAP7_75t_R%C1
cc_59 N_C1_1 N_C2_1 0.00129659f
cc_60 N_C1_4 N_C2_4 0.004121f
cc_61 N_MM9_g N_MM8_g 0.00619612f
x_PM_AOI333xp33_ASAP7_75t_R%A3 VSS A3 N_MM15_g N_A3_4 N_A3_1
+ PM_AOI333xp33_ASAP7_75t_R%A3
cc_62 N_A3_4 N_B3_1 0.000819507f
cc_63 N_MM15_g N_MM4_g 0.00327427f
cc_64 N_A3_4 N_B3_4 0.00410358f
x_PM_AOI333xp33_ASAP7_75t_R%A1 VSS A1 N_MM1_g N_A1_1 N_A1_4
+ PM_AOI333xp33_ASAP7_75t_R%A1
cc_65 N_A1_1 N_A2_1 0.00128153f
cc_66 N_A1_4 N_A2_4 0.00344193f
cc_67 N_MM1_g N_MM0_g 0.00605621f
x_PM_AOI333xp33_ASAP7_75t_R%B3 VSS B3 N_MM4_g N_B3_1 N_B3_4
+ PM_AOI333xp33_ASAP7_75t_R%B3
cc_68 N_B3_1 N_B2_1 0.0013036f
cc_69 N_B3_4 N_B2_4 0.00334931f
cc_70 N_MM4_g N_MM5_g 0.00600029f
x_PM_AOI333xp33_ASAP7_75t_R%A2 VSS A2 N_MM0_g N_A2_1 N_A2_4
+ PM_AOI333xp33_ASAP7_75t_R%A2
cc_71 N_A2_1 N_A3_1 0.00133388f
cc_72 N_A2_4 N_A3_4 0.00343854f
cc_73 N_MM0_g N_MM15_g 0.00608709f
x_PM_AOI333xp33_ASAP7_75t_R%Y VSS Y N_MM17_d N_MM12_d N_MM14_d N_MM1_d N_MM15_d
+ N_MM0_d N_Y_17 N_Y_13 N_Y_1 N_Y_18 N_Y_2 N_Y_15 N_Y_16 N_Y_4 N_Y_3 N_Y_19
+ N_Y_14 PM_AOI333xp33_ASAP7_75t_R%Y
cc_74 N_Y_17 N_MM9_g 0.000631083f
cc_75 N_Y_13 N_C1_1 0.000746162f
cc_76 N_Y_1 N_C1_4 0.00120925f
cc_77 N_Y_1 N_MM9_g 0.00153921f
cc_78 N_Y_13 N_MM9_g 0.0352028f
cc_79 N_Y_13 N_B1_1 0.000870926f
cc_80 N_Y_17 N_B1_4 0.00127474f
cc_81 N_Y_1 N_MM6_g 0.00151808f
cc_82 N_Y_1 N_B1_4 0.00169986f
cc_83 N_Y_13 N_MM6_g 0.0351116f
cc_84 N_Y_13 N_B2_4 0.000397726f
cc_85 N_Y_17 N_B2_4 0.00344617f
cc_86 N_Y_17 N_B3_4 0.00321552f
cc_87 N_Y_18 N_A3_4 0.000696609f
cc_88 N_Y_2 N_MM15_g 0.000895473f
cc_89 N_Y_17 N_A3_4 0.00138326f
cc_90 N_Y_2 N_A3_4 0.00219484f
cc_91 N_Y_15 N_MM15_g 0.0354182f
cc_92 N_Y_2 N_MM0_g 0.00128361f
cc_93 N_Y_15 N_A2_1 0.000888761f
cc_94 N_Y_18 N_A2_4 0.0011567f
cc_95 N_Y_17 N_A2_4 0.00149689f
cc_96 N_Y_2 N_A2_4 0.00267188f
cc_97 N_Y_15 N_MM0_g 0.0353181f
cc_98 N_Y_16 N_MM1_g 0.0156599f
cc_99 N_Y_4 N_A1_1 0.000919786f
cc_100 N_Y_4 N_MM1_g 0.00100932f
cc_101 N_Y_18 N_A1_4 0.00116803f
cc_102 N_Y_17 N_A1_4 0.00123243f
cc_103 N_Y_3 N_MM1_g 0.00166311f
cc_104 N_Y_16 N_A1_1 0.00174113f
cc_105 N_Y_19 N_A1_4 0.00668787f
cc_106 N_Y_14 N_MM1_g 0.05421f
cc_107 N_Y_4 N_NET030_13 0.00029755f
cc_108 N_Y_16 N_NET030_13 0.000550832f
cc_109 N_Y_15 N_NET030_11 0.00166822f
cc_110 N_Y_18 N_NET030_3 0.000701933f
cc_111 N_Y_2 N_NET030_13 0.000769361f
cc_112 N_Y_15 N_NET030_12 0.00112435f
cc_113 N_Y_4 N_NET030_3 0.00130348f
cc_114 N_Y_2 N_NET030_3 0.00304802f
cc_115 N_Y_2 N_NET030_2 0.00412705f
cc_116 N_Y_18 N_NET030_13 0.0106373f
x_PM_AOI333xp33_ASAP7_75t_R%NET030 VSS N_MM6_d N_MM5_d N_MM4_d N_MM15_s N_MM0_s
+ N_MM1_s N_NET030_1 N_NET030_10 N_NET030_11 N_NET030_2 N_NET030_12 N_NET030_3
+ N_NET030_13 PM_AOI333xp33_ASAP7_75t_R%NET030
cc_117 N_NET030_1 N_MM6_g 0.000905835f
cc_118 N_NET030_10 N_MM6_g 0.0341311f
cc_119 N_NET030_10 N_B2_1 0.000715875f
cc_120 N_NET030_1 N_MM5_g 0.000905475f
cc_121 N_NET030_10 N_MM5_g 0.0337238f
cc_122 N_NET030_11 N_B3_1 0.000550066f
cc_123 N_NET030_2 N_MM4_g 0.000950582f
cc_124 N_NET030_11 N_MM4_g 0.0340403f
cc_125 N_NET030_11 N_A3_1 0.00055804f
cc_126 N_NET030_2 N_MM15_g 0.000943863f
cc_127 N_NET030_11 N_MM15_g 0.0339875f
cc_128 N_NET030_12 N_A2_1 0.000645627f
cc_129 N_NET030_3 N_MM0_g 0.000908861f
cc_130 N_NET030_12 N_MM0_g 0.0337965f
cc_131 N_NET030_12 N_A1_1 0.00065926f
cc_132 N_NET030_3 N_MM1_g 0.000904855f
cc_133 N_NET030_12 N_MM1_g 0.0336225f
cc_134 N_NET030_1 N_NET031_13 0.000673245f
cc_135 N_NET030_13 N_NET031_3 0.000683905f
cc_136 N_NET030_10 N_NET031_11 0.00111376f
cc_137 N_NET030_10 N_NET031_12 0.00111568f
cc_138 N_NET030_2 N_NET031_3 0.0013249f
cc_139 N_NET030_1 N_NET031_3 0.00276791f
cc_140 N_NET030_1 N_NET031_2 0.00425039f
cc_141 N_NET030_13 N_NET031_13 0.0103103f
*END of AOI333xp33_ASAP7_75t_R.pxi
.ENDS
** Design:	AOI33xp33_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AOI33xp33_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AOI33xp33_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AOI33xp33_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.0327792f
.ends

.subckt PM_AOI33xp33_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.0424642f
.ends

.subckt PM_AOI33xp33_ASAP7_75t_R%NET51 VSS 2 3 1
c1 1 VSS 0.000913167f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3240 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3240 $Y2=0.0675
.ends

.subckt PM_AOI33xp33_ASAP7_75t_R%NET52 VSS 2 3 1
c1 1 VSS 0.000926019f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2700 $Y2=0.0675
.ends

.subckt PM_AOI33xp33_ASAP7_75t_R%NET53 VSS 2 3 1
c1 1 VSS 0.000929879f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_AOI33xp33_ASAP7_75t_R%NET54 VSS 2 3 1
c1 1 VSS 0.000871026f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_AOI33xp33_ASAP7_75t_R%A1 VSS 8 3 1 4
c1 1 VSS 0.00444871f
c2 3 VSS 0.0715935f
c3 4 VSS 0.0159841f
r1 9 10 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1122 $X2=0.0810 $Y2=0.1350
r2 8 9 3.32295 $w=1.3e-08 $l=1.42e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0980 $X2=0.0810 $Y2=0.1122
r3 8 4 7.52037 $w=1.3e-08 $l=3.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0980 $X2=0.0810 $Y2=0.0657
r4 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r5 1 10 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AOI33xp33_ASAP7_75t_R%B1 VSS 8 3 1 4
c1 1 VSS 0.00582229f
c2 3 VSS 0.0081952f
c3 4 VSS 0.00390878f
r1 9 10 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1207 $X2=0.2430 $Y2=0.1350
r2 8 9 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1150 $X2=0.2430 $Y2=0.1207
r3 8 4 5.30507 $w=1.3e-08 $l=2.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1150 $X2=0.2430 $Y2=0.0922
r4 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r5 1 10 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AOI33xp33_ASAP7_75t_R%B3 VSS 8 3 1 4
c1 1 VSS 0.00646379f
c2 3 VSS 0.0459896f
c3 4 VSS 0.00393227f
r1 9 10 2.50679 $w=1.3e-08 $l=1.08e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1242 $X2=0.3510 $Y2=0.1350
r2 8 9 0.524677 $w=1.3e-08 $l=2.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1220 $X2=0.3510 $Y2=0.1242
r3 8 4 6.12123 $w=1.3e-08 $l=2.63e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1220 $X2=0.3510 $Y2=0.0957
r4 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r5 1 10 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
.ends

.subckt PM_AOI33xp33_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.0419634f
.ends

.subckt PM_AOI33xp33_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.00534592f
.ends

.subckt PM_AOI33xp33_ASAP7_75t_R%A2 VSS 8 3 1 4
c1 1 VSS 0.00459247f
c2 3 VSS 0.0356094f
c3 4 VSS 0.00748784f
r1 9 10 4.72209 $w=1.3e-08 $l=2.03e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1147 $X2=0.1350 $Y2=0.1350
r2 8 9 2.73998 $w=1.3e-08 $l=1.17e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1030 $X2=0.1350 $Y2=0.1147
r3 8 4 3.90593 $w=1.3e-08 $l=1.68e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1030 $X2=0.1350 $Y2=0.0862
r4 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r5 1 10 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AOI33xp33_ASAP7_75t_R%A3 VSS 11 3 1 4
c1 1 VSS 0.00564588f
c2 3 VSS 0.0349639f
c3 4 VSS 0.00475965f
r1 11 10 0.991056 $w=1.3e-08 $l=4.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1720 $X2=0.1890 $Y2=0.1677
r2 9 10 3.20636 $w=1.3e-08 $l=1.37e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1540 $X2=0.1890 $Y2=0.1677
r3 8 9 4.4306 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1540
r4 4 8 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0980 $X2=0.1890 $Y2=0.1350
r5 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r6 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AOI33xp33_ASAP7_75t_R%B2 VSS 8 3 1 4
c1 1 VSS 0.00517469f
c2 3 VSS 0.00874533f
c3 4 VSS 0.00358833f
r1 9 10 2.50679 $w=1.3e-08 $l=1.08e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1242 $X2=0.2970 $Y2=0.1350
r2 8 9 0.524677 $w=1.3e-08 $l=2.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1220 $X2=0.2970 $Y2=0.1242
r3 8 4 6.12123 $w=1.3e-08 $l=2.63e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1220 $X2=0.2970 $Y2=0.0957
r4 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r5 1 10 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_AOI33xp33_ASAP7_75t_R%NET015 VSS 16 17 33 34 37 38 1 10 13 2 11 12 3
c1 1 VSS 0.00886758f
c2 2 VSS 0.00633071f
c3 3 VSS 0.00470427f
c4 10 VSS 0.00389846f
c5 11 VSS 0.00290764f
c6 12 VSS 0.00212652f
c7 13 VSS 0.0228223f
r1 38 36 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2160 $X2=0.1225 $Y2=0.2160
r2 1 36 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2160 $X2=0.1225 $Y2=0.2160
r3 10 1 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2160 $X2=0.1080 $Y2=0.2160
r4 37 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2160 $X2=0.0935 $Y2=0.2160
r5 34 32 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2160 $X2=0.2305 $Y2=0.2160
r6 2 32 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2160 $X2=0.2305 $Y2=0.2160
r7 11 2 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2160 $X2=0.2160 $Y2=0.2160
r8 33 11 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2160 $X2=0.2015 $Y2=0.2160
r9 1 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2160
+ $X2=0.1080 $Y2=0.2340
r10 2 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2160
+ $X2=0.2160 $Y2=0.2340
r11 29 30 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.1215 $Y2=0.2340
r12 28 30 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1215 $Y2=0.2340
r13 27 28 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r14 26 27 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r15 25 26 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1995
+ $Y=0.2340 $X2=0.1890 $Y2=0.2340
r16 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2295 $Y2=0.2340
r17 22 23 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2040
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r18 22 25 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2040
+ $Y=0.2340 $X2=0.1995 $Y2=0.2340
r19 21 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2295 $Y2=0.2340
r20 20 21 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2540
+ $Y=0.2340 $X2=0.2430 $Y2=0.2340
r21 13 18 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2855
+ $Y=0.2340 $X2=0.3240 $Y2=0.2340
r22 13 20 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2855
+ $Y=0.2340 $X2=0.2540 $Y2=0.2340
r23 3 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2160
+ $X2=0.3240 $Y2=0.2340
r24 17 15 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2160 $X2=0.3385 $Y2=0.2160
r25 3 15 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2160 $X2=0.3385 $Y2=0.2160
r26 12 3 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2160 $X2=0.3240 $Y2=0.2160
r27 16 12 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2160 $X2=0.3095 $Y2=0.2160
.ends

.subckt PM_AOI33xp33_ASAP7_75t_R%Y VSS 31 20 21 45 48 49 1 13 10 14 11 2 12 15 3
c1 1 VSS 0.00605859f
c2 2 VSS 0.00286755f
c3 3 VSS 0.00413715f
c4 10 VSS 0.00284837f
c5 11 VSS 0.00214464f
c6 12 VSS 0.00236719f
c7 13 VSS 0.0193823f
c8 14 VSS 0.00191596f
c9 15 VSS 0.00424059f
c10 16 VSS 0.00339471f
c11 17 VSS 0.00110927f
r1 48 47 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2160 $X2=0.2845 $Y2=0.2160
r2 2 47 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.2160 $X2=0.2845 $Y2=0.2160
r3 11 2 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2160 $X2=0.2700 $Y2=0.2160
r4 49 11 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2160 $X2=0.2555 $Y2=0.2160
r5 12 3 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2160 $X2=0.3760 $Y2=0.2160
r6 45 12 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2160 $X2=0.3635 $Y2=0.2160
r7 2 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2160
+ $X2=0.2700 $Y2=0.1980
r8 3 35 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2160
+ $X2=0.3780 $Y2=0.1980
r9 42 43 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1980 $X2=0.2835 $Y2=0.1980
r10 40 43 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1980 $X2=0.2835 $Y2=0.1980
r11 39 40 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3220
+ $Y=0.1980 $X2=0.2970 $Y2=0.1980
r12 38 39 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3400
+ $Y=0.1980 $X2=0.3220 $Y2=0.1980
r13 37 38 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1980 $X2=0.3400 $Y2=0.1980
r14 35 36 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.1980 $X2=0.3915 $Y2=0.1980
r15 14 35 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3645
+ $Y=0.1980 $X2=0.3780 $Y2=0.1980
r16 14 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3645
+ $Y=0.1980 $X2=0.3510 $Y2=0.1980
r17 17 34 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.1980 $X2=0.4050 $Y2=0.1765
r18 17 36 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.1980 $X2=0.3915 $Y2=0.1980
r19 33 34 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1170 $X2=0.4050 $Y2=0.1765
r20 15 32 3.50163 $w=1.45753e-08 $l=1.83e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.0575 $X2=0.4050 $Y2=0.0392
r21 15 33 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0575 $X2=0.4050 $Y2=0.1170
r22 31 32 0.637778 $w=1.8e-08 $l=6.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0330 $X2=0.4050 $Y2=0.0392
r23 31 16 0.331644 $w=1.8e-08 $l=3.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0330 $X2=0.4050 $Y2=0.0297
r24 31 30 4.24844 $w=9e-09 $l=2.71662e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.0330 $X2=0.3780 $Y2=0.0360
r25 29 30 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r26 28 29 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.0360 $X2=0.3510 $Y2=0.0360
r27 27 28 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.3240 $Y2=0.0360
r28 26 27 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2720
+ $Y=0.0360 $X2=0.2970 $Y2=0.0360
r29 25 26 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2540
+ $Y=0.0360 $X2=0.2720 $Y2=0.0360
r30 24 25 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2540 $Y2=0.0360
r31 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r32 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.2295 $Y2=0.0360
r33 13 22 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2040
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r34 1 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0675
+ $X2=0.2160 $Y2=0.0360
r35 21 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r36 1 19 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r37 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r38 20 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2015 $Y2=0.0675
.ends


*
.SUBCKT AOI33xp33_ASAP7_75t_R VSS VDD A1 A2 A3 B1 B2 B3 Y
*
* VSS VSS
* VDD VDD
* A1 A1
* A2 A2
* A3 A3
* B1 B1
* B2 B2
* B3 B3
* Y Y
*
*

MM47 N_MM47_d N_MM47_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM46 N_MM46_d N_MM46_g N_MM46_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM39 N_MM39_d N_MM39_g N_MM39_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM44 N_MM44_d N_MM44_g N_MM44_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM45 N_MM45_d N_MM38_g N_MM45_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM48 N_MM48_d N_MM37_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM31 N_MM31_d N_MM47_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM32 N_MM32_d N_MM46_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM33 N_MM33_d N_MM39_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM35 N_MM35_d N_MM44_g N_MM35_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM38 N_MM38_d N_MM38_g N_MM38_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM37 N_MM37_d N_MM37_g N_MM37_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2


*include "AOI33xp33_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AOI33xp33_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AOI33xp33_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_AOI33xp33_ASAP7_75t_R%noxref_16
cc_1 N_noxref_16_1 N_MM47_g 0.00378294f
cc_2 N_noxref_16_1 N_noxref_15_1 0.00192233f
x_PM_AOI33xp33_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_AOI33xp33_ASAP7_75t_R%noxref_15
cc_3 N_noxref_15_1 N_MM47_g 0.00186768f
x_PM_AOI33xp33_ASAP7_75t_R%NET51 VSS N_MM45_s N_MM48_d N_NET51_1
+ PM_AOI33xp33_ASAP7_75t_R%NET51
cc_4 N_NET51_1 N_MM38_g 0.017314f
cc_5 N_NET51_1 N_MM37_g 0.0172179f
x_PM_AOI33xp33_ASAP7_75t_R%NET52 VSS N_MM44_s N_MM45_d N_NET52_1
+ PM_AOI33xp33_ASAP7_75t_R%NET52
cc_6 N_NET52_1 N_MM44_g 0.0175147f
cc_7 N_NET52_1 N_MM38_g 0.0174113f
x_PM_AOI33xp33_ASAP7_75t_R%NET53 VSS N_MM47_d N_MM46_s N_NET53_1
+ PM_AOI33xp33_ASAP7_75t_R%NET53
cc_8 N_NET53_1 N_MM47_g 0.0174821f
cc_9 N_NET53_1 N_MM46_g 0.0174392f
x_PM_AOI33xp33_ASAP7_75t_R%NET54 VSS N_MM46_d N_MM39_s N_NET54_1
+ PM_AOI33xp33_ASAP7_75t_R%NET54
cc_10 N_NET54_1 N_MM46_g 0.0173889f
cc_11 N_NET54_1 N_MM39_g 0.017246f
x_PM_AOI33xp33_ASAP7_75t_R%A1 VSS A1 N_MM47_g N_A1_1 N_A1_4
+ PM_AOI33xp33_ASAP7_75t_R%A1
x_PM_AOI33xp33_ASAP7_75t_R%B1 VSS B1 N_MM44_g N_B1_1 N_B1_4
+ PM_AOI33xp33_ASAP7_75t_R%B1
cc_12 N_B1_1 N_A3_1 0.00111168f
cc_13 N_B1_4 N_A3_4 0.00379739f
cc_14 N_MM44_g N_MM39_g 0.00623789f
x_PM_AOI33xp33_ASAP7_75t_R%B3 VSS B3 N_MM37_g N_B3_1 N_B3_4
+ PM_AOI33xp33_ASAP7_75t_R%B3
cc_15 N_B3_1 N_B2_1 0.00157572f
cc_16 N_B3_4 N_B2_4 0.00370094f
cc_17 N_MM37_g N_MM38_g 0.00838822f
x_PM_AOI33xp33_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_AOI33xp33_ASAP7_75t_R%noxref_17
cc_18 N_noxref_17_1 N_MM37_g 0.00159521f
cc_19 N_noxref_17_1 N_Y_15 0.000943037f
x_PM_AOI33xp33_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_AOI33xp33_ASAP7_75t_R%noxref_18
cc_20 N_noxref_18_1 N_MM37_g 0.00346645f
cc_21 N_noxref_18_1 N_Y_12 0.0279007f
cc_22 N_noxref_18_1 N_noxref_17_1 0.00189429f
x_PM_AOI33xp33_ASAP7_75t_R%A2 VSS A2 N_MM46_g N_A2_1 N_A2_4
+ PM_AOI33xp33_ASAP7_75t_R%A2
cc_23 N_A2_1 N_MM47_g 0.00126092f
cc_24 N_A2_1 N_A1_1 0.00164722f
cc_25 N_A2_4 N_A1_4 0.00635302f
cc_26 N_MM46_g N_MM47_g 0.00731835f
x_PM_AOI33xp33_ASAP7_75t_R%A3 VSS A3 N_MM39_g N_A3_1 N_A3_4
+ PM_AOI33xp33_ASAP7_75t_R%A3
cc_27 N_A3_1 N_A2_1 0.00147811f
cc_28 N_A3_4 N_A2_4 0.00538151f
cc_29 N_MM39_g N_MM46_g 0.00842516f
x_PM_AOI33xp33_ASAP7_75t_R%B2 VSS B2 N_MM38_g N_B2_1 N_B2_4
+ PM_AOI33xp33_ASAP7_75t_R%B2
cc_30 N_B2_1 N_B1_1 0.00157088f
cc_31 N_B2_4 N_B1_4 0.00363445f
cc_32 N_MM38_g N_MM44_g 0.008316f
x_PM_AOI33xp33_ASAP7_75t_R%NET015 VSS N_MM38_s N_MM37_s N_MM33_d N_MM35_s
+ N_MM31_d N_MM32_d N_NET015_1 N_NET015_10 N_NET015_13 N_NET015_2 N_NET015_11
+ N_NET015_12 N_NET015_3 PM_AOI33xp33_ASAP7_75t_R%NET015
cc_33 N_NET015_1 N_MM47_g 0.000719083f
cc_34 N_NET015_1 N_A1_4 0.000982103f
cc_35 N_NET015_10 N_MM47_g 0.0252494f
cc_36 N_NET015_13 N_A2_4 0.00111441f
cc_37 N_NET015_1 N_A2_4 0.00150306f
cc_38 N_NET015_10 N_MM46_g 0.0254323f
cc_39 N_NET015_13 N_A3_4 0.00121917f
cc_40 N_NET015_2 N_A3_4 0.0015792f
cc_41 N_NET015_11 N_MM39_g 0.0254301f
cc_42 N_NET015_2 N_MM44_g 0.00051421f
cc_43 N_NET015_11 N_MM44_g 0.0250869f
cc_44 N_NET015_12 N_MM38_g 0.0253293f
cc_45 N_NET015_12 N_MM37_g 0.0250007f
x_PM_AOI33xp33_ASAP7_75t_R%Y VSS Y N_MM39_d N_MM44_d N_MM37_d N_MM38_d N_MM35_d
+ N_Y_1 N_Y_13 N_Y_10 N_Y_14 N_Y_11 N_Y_2 N_Y_12 N_Y_15 N_Y_3
+ PM_AOI33xp33_ASAP7_75t_R%Y
cc_46 N_Y_1 N_MM46_g 0.000338828f
cc_47 N_Y_1 N_A2_4 0.00136036f
cc_48 N_Y_13 N_A3_4 0.000598047f
cc_49 N_Y_10 N_A3_1 0.000642192f
cc_50 N_Y_1 N_A3_4 0.00146678f
cc_51 N_Y_1 N_MM39_g 0.00155917f
cc_52 N_Y_10 N_MM39_g 0.0358918f
cc_53 N_Y_1 N_B1_1 0.000472794f
cc_54 N_Y_14 N_B1_4 0.000587997f
cc_55 N_Y_10 N_B1_1 0.00108834f
cc_56 N_Y_13 N_B1_4 0.00123575f
cc_57 N_Y_1 N_MM44_g 0.00155666f
cc_58 N_Y_1 N_B1_4 0.00247187f
cc_59 N_Y_11 N_MM44_g 0.0108249f
cc_60 N_Y_10 N_MM44_g 0.0497616f
cc_61 N_Y_14 N_B2_1 0.000372382f
cc_62 N_Y_11 N_B2_1 0.000436533f
cc_63 N_Y_2 N_MM38_g 0.000452247f
cc_64 N_Y_14 N_B2_4 0.00125168f
cc_65 N_Y_13 N_B2_4 0.0041096f
cc_66 N_Y_11 N_MM38_g 0.0259591f
cc_67 N_Y_12 N_B3_1 0.000515187f
cc_68 N_Y_15 N_B3_1 0.000534211f
cc_69 N_Y_14 N_B3_4 0.00122952f
cc_70 N_Y_13 N_B3_4 0.00125309f
cc_71 N_Y_15 N_B3_4 0.00615983f
cc_72 N_Y_12 N_MM37_g 0.0257044f
cc_73 N_Y_11 N_NET015_13 0.000421404f
cc_74 N_Y_2 N_NET015_13 0.000675408f
cc_75 N_Y_11 N_NET015_11 0.000827524f
cc_76 N_Y_11 N_NET015_12 0.000846144f
cc_77 N_Y_14 N_NET015_3 0.000874146f
cc_78 N_Y_3 N_NET015_3 0.000946408f
cc_79 N_Y_2 N_NET015_3 0.00231492f
cc_80 N_Y_2 N_NET015_2 0.00310329f
cc_81 N_Y_14 N_NET015_13 0.00974594f
*END of AOI33xp33_ASAP7_75t_R.pxi
.ENDS
** Design:	A2O1A1Ixp33_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "A2O1A1Ixp33_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "A2O1A1Ixp33_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_A2O1A1Ixp33_ASAP7_75t_R%NET015 VSS 2 3 1
c1 1 VSS 0.00101967f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_A2O1A1Ixp33_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.00602328f
.ends

.subckt PM_A2O1A1Ixp33_ASAP7_75t_R%A1 VSS 9 3 1 4
c1 1 VSS 0.00269054f
c2 3 VSS 0.0432751f
c3 4 VSS 0.0147614f
r1 9 8 1.92382 $w=1.3e-08 $l=8.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1600 $X2=0.0810 $Y2=0.1517
r2 7 8 3.90593 $w=1.3e-08 $l=1.67e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1517
r3 4 7 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0980 $X2=0.0810 $Y2=0.1350
r4 6 7 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1355
+ $X2=0.0810 $Y2=0.1350
r5 3 1 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1 $thickness=5.5619e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0810 $Y2=0.1245
r6 1 6 6.49795 $w=1.53e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08 $X=0.0810
+ $Y=0.1245 $X2=0.0810 $Y2=0.1355
.ends

.subckt PM_A2O1A1Ixp33_ASAP7_75t_R%A2 VSS 9 3 1 4
c1 1 VSS 0.00719274f
c2 3 VSS 0.0832909f
c3 4 VSS 0.00486209f
r1 9 8 0.874462 $w=1.3e-08 $l=3.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1520 $X2=0.1350 $Y2=0.1482
r2 7 8 2.85657 $w=1.3e-08 $l=1.22e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1360 $X2=0.1350 $Y2=0.1482
r3 4 7 8.74462 $w=1.3e-08 $l=3.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0985 $X2=0.1350 $Y2=0.1360
r4 3 1 6.51726 $w=1.18568e-07 $l=5e-10 $layer=LIG $thickness=5.19024e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1350 $Y2=0.1355
r5 1 7 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1355
+ $X2=0.1350 $Y2=0.1360
.ends

.subckt PM_A2O1A1Ixp33_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.00603763f
.ends

.subckt PM_A2O1A1Ixp33_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.0316034f
.ends

.subckt PM_A2O1A1Ixp33_ASAP7_75t_R%B VSS 6 3 4 1
c1 1 VSS 0.0089266f
c2 3 VSS 0.0459767f
c3 4 VSS 0.00561697f
r1 7 8 3.08976 $w=1.3e-08 $l=1.33e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1227 $X2=0.1890 $Y2=0.1360
r2 6 7 1.10765 $w=1.3e-08 $l=4.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1180 $X2=0.1890 $Y2=0.1227
r3 6 4 4.37231 $w=1.3e-08 $l=1.88e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1180 $X2=0.1890 $Y2=0.0992
r4 3 1 6.81262 $w=1.1611e-07 $l=1e-09 $layer=LIG $thickness=5.18095e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1890 $Y2=0.1360
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1360
+ $X2=0.1890 $Y2=0.1360
.ends

.subckt PM_A2O1A1Ixp33_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00484912f
.ends

.subckt PM_A2O1A1Ixp33_ASAP7_75t_R%NET06 VSS 11 25 28 7 9 1 2 8
c1 1 VSS 0.00639396f
c2 2 VSS 0.00715135f
c3 7 VSS 0.00312007f
c4 8 VSS 0.00330288f
c5 9 VSS 0.0187564f
r1 28 27 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r2 26 27 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2260 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r3 2 26 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2140 $Y=0.0675 $X2=0.2260 $Y2=0.0675
r4 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0675 $X2=0.2140 $Y2=0.0675
r5 25 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2015 $Y2=0.0675
r6 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0675
+ $X2=0.2195 $Y2=0.0360
r7 21 22 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2105
+ $Y=0.0360 $X2=0.2195 $Y2=0.0360
r8 20 21 1.86552 $w=1.3e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.2025
+ $Y=0.0360 $X2=0.2105 $Y2=0.0360
r9 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.2025 $Y2=0.0360
r10 18 19 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1780
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r11 17 18 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1600
+ $Y=0.0360 $X2=0.1780 $Y2=0.0360
r12 16 17 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1600 $Y2=0.0360
r13 15 16 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r14 14 15 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0360 $X2=0.1080 $Y2=0.0360
r15 13 14 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0675
+ $Y=0.0360 $X2=0.0810 $Y2=0.0360
r16 12 13 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.0360 $X2=0.0675 $Y2=0.0360
r17 9 12 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r18 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0540 $Y2=0.0360
r19 11 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r20 7 10 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r21 1 7 1e-05
.ends

.subckt PM_A2O1A1Ixp33_ASAP7_75t_R%Y VSS 22 16 34 37 8 1 9 11 2 12 7 13
c1 1 VSS 0.00999012f
c2 2 VSS 0.0052336f
c3 7 VSS 0.0021394f
c4 8 VSS 0.00203141f
c5 9 VSS 0.00039238f
c6 10 VSS 2.32571e-20
c7 11 VSS 0.00541036f
c8 12 VSS 0.00334268f
c9 13 VSS 0.00382422f
c10 14 VSS 0.00253643f
r1 39 40 0.264706 $w=1.7e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2260 $Y=0.1975 $X2=0.2305 $Y2=0.1975
r2 1 39 0.705882 $w=1.7e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2140 $Y=0.1975 $X2=0.2260 $Y2=0.1975
r3 10 1 0.735294 $w=1.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.1975 $X2=0.2140 $Y2=0.1975
r4 37 36 0.0675676 $w=3.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2245 $X2=0.2305 $Y2=0.2245
r5 1 36 0.391892 $w=3.7e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2245 $X2=0.2305 $Y2=0.2245
r6 1 40 0.471383 $w=3.35517e-08 $l=3.06472e-08 $layer=P_src_drn
+ $thickness=1e-09 $X=0.2160 $Y=0.2245 $X2=0.2305 $Y2=0.1975
r7 9 1 0.391892 $w=3.7e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2245 $X2=0.2160 $Y2=0.2245
r8 8 1 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.1755 $X2=0.2140 $Y2=0.1755
r9 34 8 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.1755 $X2=0.2015 $Y2=0.1755
r10 1 31 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2220 $Y=0.2160
+ $X2=0.2245 $Y2=0.2240
r11 29 31 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2320
+ $Y=0.2240 $X2=0.2245 $Y2=0.2240
r12 27 28 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2355
+ $Y=0.2240 $X2=0.2445 $Y2=0.2240
r13 27 29 0.816164 $w=1.3e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2355
+ $Y=0.2240 $X2=0.2320 $Y2=0.2240
r14 26 28 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2570
+ $Y=0.2240 $X2=0.2445 $Y2=0.2240
r15 11 14 3.48106 $w=1.50455e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2750 $Y=0.2240 $X2=0.2970 $Y2=0.2240
r16 11 26 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2750
+ $Y=0.2240 $X2=0.2570 $Y2=0.2240
r17 14 25 2.19852 $w=1.83455e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.2240 $X2=0.2970 $Y2=0.2075
r18 24 25 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1950 $X2=0.2970 $Y2=0.2075
r19 23 24 2.62338 $w=1.3e-08 $l=1.13e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1837 $X2=0.2970 $Y2=0.1950
r20 22 23 1.57403 $w=1.3e-08 $l=6.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1770 $X2=0.2970 $Y2=0.1837
r21 22 21 11.2514 $w=1.3e-08 $l=4.83e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1770 $X2=0.2970 $Y2=0.1287
r22 20 21 12.4174 $w=1.3e-08 $l=5.32e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0755 $X2=0.2970 $Y2=0.1287
r23 12 19 2.66732 $w=1.57273e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0625 $X2=0.2970 $Y2=0.0460
r24 12 20 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0625 $X2=0.2970 $Y2=0.0755
r25 18 19 1.26818 $w=1.72857e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2865 $Y=0.0460 $X2=0.2970 $Y2=0.0460
r26 17 18 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2760
+ $Y=0.0460 $X2=0.2865 $Y2=0.0460
r27 13 17 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2645
+ $Y=0.0460 $X2=0.2760 $Y2=0.0460
r28 2 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2730 $Y=0.0675
+ $X2=0.2760 $Y2=0.0460
r29 7 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2680 $Y2=0.0675
r30 16 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
.ends

.subckt PM_A2O1A1Ixp33_ASAP7_75t_R%C VSS 6 3 4 1
c1 1 VSS 0.00692623f
c2 3 VSS 0.0346322f
c3 4 VSS 0.00471362f
r1 7 8 7.17059 $w=1.3e-08 $l=3.08e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1052 $X2=0.2430 $Y2=0.1360
r2 6 7 5.18847 $w=1.3e-08 $l=2.22e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0830 $X2=0.2430 $Y2=0.1052
r3 6 4 0.291487 $w=1.3e-08 $l=1.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0830 $X2=0.2430 $Y2=0.0817
r4 3 1 6.81262 $w=1.1611e-07 $l=1e-09 $layer=LIG $thickness=5.18095e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2430 $Y2=0.1360
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1360
+ $X2=0.2430 $Y2=0.1360
.ends

.subckt PM_A2O1A1Ixp33_ASAP7_75t_R%NET2 VSS 11 22 23 7 9 1 2 8
c1 1 VSS 0.00846087f
c2 2 VSS 0.00750698f
c3 7 VSS 0.00395737f
c4 8 VSS 0.00344709f
c5 9 VSS 0.0135525f
r1 23 21 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r2 2 21 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r4 22 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r5 2 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r6 17 18 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r7 16 17 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1485 $Y2=0.2340
r8 15 16 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r9 14 15 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.2340 $X2=0.1080 $Y2=0.2340
r10 13 14 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0675
+ $Y=0.2340 $X2=0.0810 $Y2=0.2340
r11 12 13 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2340 $X2=0.0675 $Y2=0.2340
r12 9 12 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r13 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r14 11 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r15 7 10 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r16 1 7 1e-05
.ends


*
.SUBCKT A2O1A1Ixp33_ASAP7_75t_R VSS VDD A1 A2 B C Y
*
* VSS VSS
* VDD VDD
* A1 A1
* A2 A2
* B B
* C C
* Y Y
*
*

MM0 N_MM0_d N_MM0_g N_MM0_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM1_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM7_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2


*include "A2O1A1Ixp33_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "A2O1A1Ixp33_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_A2O1A1Ixp33_ASAP7_75t_R%NET015 VSS N_MM0_s N_MM1_d N_NET015_1
+ PM_A2O1A1Ixp33_ASAP7_75t_R%NET015
cc_1 N_NET015_1 N_MM0_g 0.0172765f
cc_2 N_NET015_1 N_MM1_g 0.0171858f
x_PM_A2O1A1Ixp33_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_A2O1A1Ixp33_ASAP7_75t_R%noxref_12
cc_3 N_noxref_12_1 N_MM0_g 0.00162707f
cc_4 N_noxref_12_1 N_NET06_7 0.000560257f
cc_5 N_noxref_12_1 N_NET2_7 0.0363526f
cc_6 N_noxref_12_1 N_noxref_11_1 0.00179454f
x_PM_A2O1A1Ixp33_ASAP7_75t_R%A1 VSS A1 N_MM0_g N_A1_1 N_A1_4
+ PM_A2O1A1Ixp33_ASAP7_75t_R%A1
x_PM_A2O1A1Ixp33_ASAP7_75t_R%A2 VSS A2 N_MM1_g N_A2_1 N_A2_4
+ PM_A2O1A1Ixp33_ASAP7_75t_R%A2
cc_7 N_A2_1 N_A1_1 0.00122161f
cc_8 N_A2_4 N_A1_4 0.00483287f
cc_9 N_MM1_g N_MM0_g 0.00603323f
x_PM_A2O1A1Ixp33_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_A2O1A1Ixp33_ASAP7_75t_R%noxref_11
cc_10 N_noxref_11_1 N_MM0_g 0.00163126f
cc_11 N_noxref_11_1 N_NET06_7 0.0363284f
cc_12 N_noxref_11_1 N_NET2_7 0.000563921f
x_PM_A2O1A1Ixp33_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_A2O1A1Ixp33_ASAP7_75t_R%noxref_14
cc_13 N_noxref_14_1 N_MM2_g 0.00341634f
cc_14 N_noxref_14_1 N_Y_9 0.00165522f
cc_15 N_noxref_14_1 N_noxref_13_1 0.00189001f
x_PM_A2O1A1Ixp33_ASAP7_75t_R%B VSS B N_MM7_g N_B_4 N_B_1
+ PM_A2O1A1Ixp33_ASAP7_75t_R%B
cc_16 N_MM7_g N_MM1_g 0.00326146f
cc_17 N_B_4 N_A2_4 0.00612064f
x_PM_A2O1A1Ixp33_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_A2O1A1Ixp33_ASAP7_75t_R%noxref_13
cc_18 N_noxref_13_1 N_MM2_g 0.00157696f
cc_19 N_noxref_13_1 N_Y_2 0.000940452f
cc_20 N_noxref_13_1 N_Y_7 0.0373049f
x_PM_A2O1A1Ixp33_ASAP7_75t_R%NET06 VSS N_MM0_d N_MM7_d N_MM2_s N_NET06_7
+ N_NET06_9 N_NET06_1 N_NET06_2 N_NET06_8 PM_A2O1A1Ixp33_ASAP7_75t_R%NET06
cc_21 N_NET06_7 N_A1_1 0.000930519f
cc_22 N_NET06_9 N_A1_4 0.00134336f
cc_23 N_NET06_1 N_MM0_g 0.00180903f
cc_24 N_NET06_1 N_A1_4 0.00220011f
cc_25 N_NET06_7 N_MM0_g 0.0348993f
cc_26 N_NET06_9 N_A2_4 0.00358262f
cc_27 N_NET06_9 N_B_4 0.00112831f
cc_28 N_NET06_2 N_MM7_g 0.00114094f
cc_29 N_NET06_2 N_B_4 0.00159954f
cc_30 N_NET06_8 N_MM7_g 0.0346539f
cc_31 N_NET06_2 N_C_4 0.000776797f
cc_32 N_NET06_2 N_MM2_g 0.00107091f
cc_33 N_NET06_8 N_MM2_g 0.0346408f
x_PM_A2O1A1Ixp33_ASAP7_75t_R%Y VSS Y N_MM2_d N_MM5_d N_MM6_d N_Y_8 N_Y_1 N_Y_9
+ N_Y_11 N_Y_2 N_Y_12 N_Y_7 N_Y_13 PM_A2O1A1Ixp33_ASAP7_75t_R%Y
cc_34 N_Y_8 N_B_1 0.00081978f
cc_35 N_Y_1 N_B_4 0.00124543f
cc_36 N_Y_1 N_MM7_g 0.00126526f
cc_37 N_Y_8 N_MM7_g 0.00966043f
cc_38 N_Y_9 N_MM7_g 0.0253719f
cc_39 N_Y_1 N_C_1 0.00273745f
cc_40 N_Y_11 N_C_4 0.00092629f
cc_41 N_Y_2 N_MM2_g 0.00127339f
cc_42 N_Y_1 N_MM2_g 0.00228664f
cc_43 N_Y_9 N_MM2_g 0.00519046f
cc_44 N_Y_12 N_C_4 0.00712807f
cc_45 N_Y_8 N_MM2_g 0.0099723f
cc_46 N_Y_7 N_MM2_g 0.0552396f
cc_47 N_Y_7 N_NET06_8 0.000607176f
cc_48 N_Y_13 N_NET06_9 0.00101479f
cc_49 N_Y_2 N_NET06_8 0.00133913f
cc_50 N_Y_2 N_NET06_2 0.00278244f
cc_51 N_Y_11 N_NET2_9 0.000688379f
cc_52 N_Y_1 N_NET2_2 0.00123757f
cc_53 N_Y_1 N_NET2_8 0.00296962f
x_PM_A2O1A1Ixp33_ASAP7_75t_R%C VSS C N_MM2_g N_C_4 N_C_1
+ PM_A2O1A1Ixp33_ASAP7_75t_R%C
cc_54 N_MM2_g N_MM7_g 0.0032594f
cc_55 N_C_4 N_B_4 0.00575622f
x_PM_A2O1A1Ixp33_ASAP7_75t_R%NET2 VSS N_MM3_d N_MM4_d N_MM5_s N_NET2_7 N_NET2_9
+ N_NET2_1 N_NET2_2 N_NET2_8 PM_A2O1A1Ixp33_ASAP7_75t_R%NET2
cc_56 N_NET2_7 N_A1_1 0.000658108f
cc_57 N_NET2_9 N_A1_4 0.00127906f
cc_58 N_NET2_1 N_MM0_g 0.0014901f
cc_59 N_NET2_1 N_A1_4 0.00195371f
cc_60 N_NET2_7 N_MM0_g 0.0343766f
cc_61 N_NET2_9 N_A2_4 0.00112377f
cc_62 N_NET2_2 N_MM1_g 0.00119998f
cc_63 N_NET2_2 N_A2_4 0.00158558f
cc_64 N_NET2_8 N_MM1_g 0.0347537f
cc_65 N_NET2_8 N_B_1 0.00078495f
cc_66 N_NET2_2 N_B_4 0.00100968f
cc_67 N_NET2_2 N_MM7_g 0.00119672f
cc_68 N_NET2_8 N_MM7_g 0.0344607f
*END of A2O1A1Ixp33_ASAP7_75t_R.pxi
.ENDS
** Design:	A2O1A1O1Ixp25_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "A2O1A1O1Ixp25_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "A2O1A1O1Ixp25_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_A2O1A1O1Ixp25_ASAP7_75t_R%NET25 VSS 2 3 1
c1 1 VSS 0.0010007f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_A2O1A1O1Ixp25_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.0423347f
.ends

.subckt PM_A2O1A1O1Ixp25_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00607742f
.ends

.subckt PM_A2O1A1O1Ixp25_ASAP7_75t_R%A1 VSS 8 3 1 4
c1 1 VSS 0.00729957f
c2 3 VSS 0.0833026f
c3 4 VSS 0.00510021f
r1 8 7 5.18847 $w=1.3e-08 $l=2.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1880 $X2=0.1350 $Y2=0.1657
r2 6 7 7.17059 $w=1.3e-08 $l=3.07e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1657
r3 4 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0980 $X2=0.1350 $Y2=0.1350
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r5 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_A2O1A1O1Ixp25_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00599161f
.ends

.subckt PM_A2O1A1O1Ixp25_ASAP7_75t_R%A2 VSS 6 3 1 4
c1 1 VSS 0.00309665f
c2 3 VSS 0.0432855f
c3 4 VSS 0.0149888f
r1 7 8 7.17059 $w=1.3e-08 $l=3.08e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1042 $X2=0.0810 $Y2=0.1350
r2 6 7 5.18847 $w=1.3e-08 $l=2.22e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0820 $X2=0.0810 $Y2=0.1042
r3 6 4 1.45744 $w=1.3e-08 $l=6.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0820 $X2=0.0810 $Y2=0.0757
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_A2O1A1O1Ixp25_ASAP7_75t_R%NET4 VSS 11 21 22 7 9 1 2 8
c1 1 VSS 0.00842285f
c2 2 VSS 0.00757815f
c3 7 VSS 0.00396938f
c4 8 VSS 0.00339874f
c5 9 VSS 0.0126378f
r1 22 20 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r2 2 20 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r4 21 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r5 2 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r6 17 18 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r7 16 17 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1485 $Y2=0.2340
r8 15 16 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r9 14 15 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.2340 $X2=0.1080 $Y2=0.2340
r10 13 14 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0675
+ $Y=0.2340 $X2=0.0810 $Y2=0.2340
r11 12 13 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2340 $X2=0.0675 $Y2=0.2340
r12 9 12 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r13 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r14 11 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r15 7 10 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r16 1 7 1e-05
.ends

.subckt PM_A2O1A1O1Ixp25_ASAP7_75t_R%B VSS 8 3 4
c1 1 VSS 0.0091262f
c2 3 VSS 0.0460281f
c3 4 VSS 0.00595106f
r1 8 7 1.22425 $w=1.3e-08 $l=5.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1540 $X2=0.1890 $Y2=0.1487
r2 6 7 3.20636 $w=1.3e-08 $l=1.37e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1487
r3 4 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0980 $X2=0.1890 $Y2=0.1350
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r5 1 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_A2O1A1O1Ixp25_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00569283f
.ends

.subckt PM_A2O1A1O1Ixp25_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.00538645f
.ends

.subckt PM_A2O1A1O1Ixp25_ASAP7_75t_R%D VSS 7 3 1 5 6 4
c1 1 VSS 0.00604647f
c2 3 VSS 0.0445743f
c3 4 VSS 0.00319363f
c4 5 VSS 0.00328278f
c5 6 VSS 0.00261915f
c6 7 VSS 0.00319569f
r1 7 5 7.33112 $w=1.42329e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.1360 $X2=0.3510 $Y2=0.1725
r2 7 4 7.56431 $w=1.42e-08 $l=3.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1360 $X2=0.3510 $Y2=0.0985
r3 7 12 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1360 $X2=0.3735 $Y2=0.1360
r4 6 11 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3915
+ $Y=0.1360 $X2=0.4050 $Y2=0.1360
r5 6 12 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3915
+ $Y=0.1360 $X2=0.3735 $Y2=0.1360
r6 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r7 1 11 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1360
.ends

.subckt PM_A2O1A1O1Ixp25_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.0418935f
.ends

.subckt PM_A2O1A1O1Ixp25_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.00551495f
.ends

.subckt PM_A2O1A1O1Ixp25_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.00662321f
.ends

.subckt PM_A2O1A1O1Ixp25_ASAP7_75t_R%NET12 VSS 11 24 25 7 9 1 2 8
c1 1 VSS 0.00644995f
c2 2 VSS 0.00731365f
c3 7 VSS 0.00313513f
c4 8 VSS 0.00345892f
c5 9 VSS 0.0183145f
r1 25 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r2 2 23 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r4 24 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2015 $Y2=0.0675
r5 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0675
+ $X2=0.2160 $Y2=0.0360
r6 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2025
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r7 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.2025 $Y2=0.0360
r8 18 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1755
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r9 17 18 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1575
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r10 16 17 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1575 $Y2=0.0360
r11 15 16 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r12 14 15 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0360 $X2=0.1080 $Y2=0.0360
r13 13 14 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0675
+ $Y=0.0360 $X2=0.0810 $Y2=0.0360
r14 12 13 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.0360 $X2=0.0675 $Y2=0.0360
r15 9 12 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r16 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0540 $Y2=0.0360
r17 11 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r18 7 10 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r19 1 7 1e-05
.ends

.subckt PM_A2O1A1O1Ixp25_ASAP7_75t_R%NET15 VSS 12 13 22 1 7 9 8 2
c1 1 VSS 0.00723819f
c2 2 VSS 0.00527212f
c3 7 VSS 0.00351688f
c4 8 VSS 0.0026575f
c5 9 VSS 0.0168228f
r1 22 21 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r2 8 21 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3800 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r3 2 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.2340
r4 19 20 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3645
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r5 18 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.2340 $X2=0.3645 $Y2=0.2340
r6 17 18 11.5429 $w=1.3e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.3015
+ $Y=0.2340 $X2=0.3510 $Y2=0.2340
r7 16 17 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.2340 $X2=0.3015 $Y2=0.2340
r8 15 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2565 $Y2=0.2340
r9 14 15 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.2340 $X2=0.2430 $Y2=0.2340
r10 9 14 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2295 $Y2=0.2340
r11 1 9 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.2340
r12 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r13 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r14 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r15 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r16 2 8 1e-05
.ends

.subckt PM_A2O1A1O1Ixp25_ASAP7_75t_R%Y VSS 26 18 28 37 13 10 1 12 2 3 14 11 15
c1 1 VSS 0.00583501f
c2 2 VSS 0.00772398f
c3 3 VSS 0.00559363f
c4 10 VSS 0.0029509f
c5 11 VSS 0.00354043f
c6 12 VSS 0.00256258f
c7 13 VSS 0.0180804f
c8 14 VSS 0.00524264f
c9 15 VSS 0.00558882f
c10 16 VSS 0.00353698f
r1 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4300 $Y2=0.2025
r2 37 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r3 3 34 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.2340
r4 34 35 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4455 $Y2=0.2340
r5 15 33 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.2340 $X2=0.4590 $Y2=0.2125
r6 15 35 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.2340 $X2=0.4455 $Y2=0.2340
r7 32 33 9.32759 $w=1.3e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1725 $X2=0.4590 $Y2=0.2125
r8 31 32 8.51143 $w=1.3e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1360 $X2=0.4590 $Y2=0.1725
r9 30 31 8.74462 $w=1.3e-08 $l=3.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0985 $X2=0.4590 $Y2=0.1360
r10 29 30 9.50248 $w=1.3e-08 $l=4.08e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0577 $X2=0.4590 $Y2=0.0985
r11 14 29 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0452 $X2=0.4590 $Y2=0.0577
r12 26 14 0.0838085 $w=1.55e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0447 $X2=0.4590 $Y2=0.0452
r13 28 27 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r14 11 27 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3800 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r15 26 16 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0447 $X2=0.4590 $Y2=0.0357
r16 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.0675
+ $X2=0.3780 $Y2=0.0360
r17 26 25 3.17357 $w=8e-09 $l=2.41234e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0447 $X2=0.4365 $Y2=0.0360
r18 24 25 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4185
+ $Y=0.0360 $X2=0.4365 $Y2=0.0360
r19 23 24 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4005
+ $Y=0.0360 $X2=0.4185 $Y2=0.0360
r20 22 23 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0360 $X2=0.4005 $Y2=0.0360
r21 21 22 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3645
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r22 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0360 $X2=0.3645 $Y2=0.0360
r23 19 20 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.3105
+ $Y=0.0360 $X2=0.3510 $Y2=0.0360
r24 13 19 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.3105 $Y2=0.0360
r25 1 13 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2700 $Y2=0.0360
r26 10 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2680 $Y2=0.0675
r27 18 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
r28 2 11 1e-05
.ends

.subckt PM_A2O1A1O1Ixp25_ASAP7_75t_R%C VSS 6 3 1 4
c1 1 VSS 0.00930852f
c2 3 VSS 0.0460871f
c3 4 VSS 0.00752999f
r1 7 8 2.85657 $w=1.3e-08 $l=1.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1227 $X2=0.2430 $Y2=0.1350
r2 6 7 0.874462 $w=1.3e-08 $l=3.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1190 $X2=0.2430 $Y2=0.1227
r3 6 4 5.77145 $w=1.3e-08 $l=2.48e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1190 $X2=0.2430 $Y2=0.0942
r4 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r5 1 8 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends


*
.SUBCKT A2O1A1O1Ixp25_ASAP7_75t_R VSS VDD A2 A1 B C D Y
*
* VSS VSS
* VDD VDD
* A2 A2
* A1 A1
* B B
* C C
* D D
* Y Y
*
*

MM1 N_MM1_d N_MM1_g N_MM1_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 VSS N_MM0_g N_MM0_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g N_MM3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM1_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM2_g N_MM7_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM4_g N_MM9_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "A2O1A1O1Ixp25_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "A2O1A1O1Ixp25_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_A2O1A1O1Ixp25_ASAP7_75t_R%NET25 VSS N_MM1_d N_MM0_s N_NET25_1
+ PM_A2O1A1O1Ixp25_ASAP7_75t_R%NET25
cc_1 N_NET25_1 N_MM1_g 0.0173468f
cc_2 N_NET25_1 N_MM0_g 0.0174531f
x_PM_A2O1A1O1Ixp25_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_A2O1A1O1Ixp25_ASAP7_75t_R%noxref_16
cc_3 N_noxref_16_1 N_MM3_g 0.00140715f
cc_4 N_noxref_16_1 N_NET15_7 0.000702209f
cc_5 N_noxref_16_1 N_noxref_15_1 0.00123759f
x_PM_A2O1A1O1Ixp25_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_A2O1A1O1Ixp25_ASAP7_75t_R%noxref_14
cc_6 N_noxref_14_1 N_MM1_g 0.00164356f
cc_7 N_noxref_14_1 N_NET12_7 0.000562511f
cc_8 N_noxref_14_1 N_NET4_7 0.0362905f
cc_9 N_noxref_14_1 N_noxref_13_1 0.00179315f
x_PM_A2O1A1O1Ixp25_ASAP7_75t_R%A1 VSS A1 N_MM0_g N_A1_1 N_A1_4
+ PM_A2O1A1O1Ixp25_ASAP7_75t_R%A1
cc_10 N_A1_1 N_A2_1 0.00130034f
cc_11 N_MM0_g N_MM1_g 0.00494269f
cc_12 N_A1_4 N_A2_4 0.006017f
x_PM_A2O1A1O1Ixp25_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_A2O1A1O1Ixp25_ASAP7_75t_R%noxref_13
cc_13 N_noxref_13_1 N_MM1_g 0.00164433f
cc_14 N_noxref_13_1 N_NET12_7 0.0364016f
cc_15 N_noxref_13_1 N_NET4_7 0.00055773f
x_PM_A2O1A1O1Ixp25_ASAP7_75t_R%A2 VSS A2 N_MM1_g N_A2_1 N_A2_4
+ PM_A2O1A1O1Ixp25_ASAP7_75t_R%A2
x_PM_A2O1A1O1Ixp25_ASAP7_75t_R%NET4 VSS N_MM6_d N_MM5_d N_MM7_s N_NET4_7
+ N_NET4_9 N_NET4_1 N_NET4_2 N_NET4_8 PM_A2O1A1O1Ixp25_ASAP7_75t_R%NET4
cc_16 N_NET4_7 N_A2_1 0.000767511f
cc_17 N_NET4_9 N_A2_4 0.00126285f
cc_18 N_NET4_1 N_MM1_g 0.00150253f
cc_19 N_NET4_1 N_A2_4 0.00213318f
cc_20 N_NET4_7 N_MM1_g 0.0343155f
cc_21 N_NET4_9 N_A1_4 0.00107857f
cc_22 N_NET4_2 N_MM0_g 0.0011785f
cc_23 N_NET4_2 N_A1_4 0.00158887f
cc_24 N_NET4_8 N_MM0_g 0.0346615f
cc_25 N_NET4_2 N_B_4 0.000944827f
cc_26 N_NET4_2 N_MM2_g 0.00117579f
cc_27 N_NET4_8 N_MM2_g 0.0350063f
x_PM_A2O1A1O1Ixp25_ASAP7_75t_R%B VSS B N_MM2_g N_B_4
+ PM_A2O1A1O1Ixp25_ASAP7_75t_R%B
cc_28 N_MM2_g N_MM0_g 0.00330438f
cc_29 N_B_4 N_A1_4 0.00627943f
x_PM_A2O1A1O1Ixp25_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_A2O1A1O1Ixp25_ASAP7_75t_R%noxref_15
cc_30 N_noxref_15_1 N_MM3_g 0.00140297f
cc_31 N_noxref_15_1 N_Y_10 0.03741f
x_PM_A2O1A1O1Ixp25_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_A2O1A1O1Ixp25_ASAP7_75t_R%noxref_20
cc_32 N_noxref_20_1 N_MM4_g 0.0014408f
cc_33 N_noxref_20_1 N_Y_12 0.0378173f
cc_34 N_noxref_20_1 N_noxref_19_1 0.00176565f
x_PM_A2O1A1O1Ixp25_ASAP7_75t_R%D VSS D N_MM4_g N_D_1 N_D_5 N_D_6 N_D_4
+ PM_A2O1A1O1Ixp25_ASAP7_75t_R%D
x_PM_A2O1A1O1Ixp25_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_A2O1A1O1Ixp25_ASAP7_75t_R%noxref_19
cc_35 N_noxref_19_1 N_MM4_g 0.0014446f
cc_36 N_noxref_19_1 N_Y_11 0.00132555f
x_PM_A2O1A1O1Ixp25_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_A2O1A1O1Ixp25_ASAP7_75t_R%noxref_17
cc_37 N_noxref_17_1 N_MM4_g 0.00159664f
cc_38 N_noxref_17_1 N_Y_11 0.0374139f
cc_39 N_noxref_17_1 N_noxref_15_1 0.00765213f
x_PM_A2O1A1O1Ixp25_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_A2O1A1O1Ixp25_ASAP7_75t_R%noxref_18
cc_40 N_noxref_18_1 N_MM4_g 0.00160107f
cc_41 N_noxref_18_1 N_NET15_8 0.0357412f
cc_42 N_noxref_18_1 N_Y_12 0.000541569f
cc_43 N_noxref_18_1 N_noxref_16_1 0.00766875f
cc_44 N_noxref_18_1 N_noxref_17_1 0.0012332f
x_PM_A2O1A1O1Ixp25_ASAP7_75t_R%NET12 VSS N_MM1_s N_MM2_d N_MM3_s N_NET12_7
+ N_NET12_9 N_NET12_1 N_NET12_2 N_NET12_8 PM_A2O1A1O1Ixp25_ASAP7_75t_R%NET12
cc_45 N_NET12_7 N_A2_1 0.000945189f
cc_46 N_NET12_9 N_A2_4 0.00138155f
cc_47 N_NET12_1 N_MM1_g 0.00182989f
cc_48 N_NET12_1 N_A2_4 0.00210531f
cc_49 N_NET12_7 N_MM1_g 0.0349992f
cc_50 N_NET12_9 N_A1_4 0.00351837f
cc_51 N_NET12_9 N_B_4 0.00113026f
cc_52 N_NET12_2 N_MM2_g 0.00116003f
cc_53 N_NET12_2 N_B_4 0.00156923f
cc_54 N_NET12_8 N_MM2_g 0.0347523f
cc_55 N_NET12_8 N_C_1 0.000663349f
cc_56 N_NET12_2 N_C_4 0.000995147f
cc_57 N_NET12_2 N_MM3_g 0.00117751f
cc_58 N_NET12_8 N_MM3_g 0.0344368f
x_PM_A2O1A1O1Ixp25_ASAP7_75t_R%NET15 VSS N_MM7_d N_MM8_d N_MM9_s N_NET15_1
+ N_NET15_7 N_NET15_9 N_NET15_8 N_NET15_2 PM_A2O1A1O1Ixp25_ASAP7_75t_R%NET15
cc_59 N_NET15_1 N_B_4 0.000957289f
cc_60 N_NET15_1 N_MM2_g 0.00116634f
cc_61 N_NET15_7 N_MM2_g 0.0348666f
cc_62 N_NET15_7 N_C_1 0.00077792f
cc_63 N_NET15_1 N_MM3_g 0.00117265f
cc_64 N_NET15_9 N_C_4 0.00131186f
cc_65 N_NET15_1 N_C_4 0.00177264f
cc_66 N_NET15_7 N_MM3_g 0.0339408f
cc_67 N_NET15_8 N_D_1 0.000714912f
cc_68 N_NET15_2 N_MM4_g 0.00171255f
cc_69 N_NET15_9 N_D_5 0.0033122f
cc_70 N_NET15_8 N_MM4_g 0.0347545f
cc_71 N_NET15_9 N_NET4_9 0.000651072f
cc_72 N_NET15_1 N_NET4_2 0.0044022f
x_PM_A2O1A1O1Ixp25_ASAP7_75t_R%Y VSS Y N_MM3_d N_MM4_d N_MM9_d N_Y_13 N_Y_10
+ N_Y_1 N_Y_12 N_Y_2 N_Y_3 N_Y_14 N_Y_11 N_Y_15 PM_A2O1A1O1Ixp25_ASAP7_75t_R%Y
cc_73 N_Y_13 N_C_4 0.000661538f
cc_74 N_Y_10 N_C_1 0.000779697f
cc_75 N_Y_1 N_C_4 0.00145564f
cc_76 N_Y_1 N_MM3_g 0.00147536f
cc_77 N_Y_10 N_MM3_g 0.0352062f
cc_78 N_Y_12 N_MM4_g 0.0156284f
cc_79 N_Y_2 N_D_5 0.000477446f
cc_80 N_Y_3 N_D_1 0.00106167f
cc_81 N_Y_3 N_MM4_g 0.00115622f
cc_82 N_Y_2 N_D_6 0.00142685f
cc_83 N_Y_12 N_D_1 0.00166324f
cc_84 N_Y_2 N_MM4_g 0.00173885f
cc_85 N_Y_13 N_D_4 0.00176882f
cc_86 N_Y_14 N_D_6 0.00183986f
cc_87 N_Y_2 N_D_4 0.00247174f
cc_88 N_Y_11 N_MM4_g 0.0547312f
cc_89 N_Y_13 N_NET12_9 0.000743838f
cc_90 N_Y_1 N_NET12_2 0.00453182f
cc_91 N_Y_12 N_NET15_8 0.000671067f
cc_92 N_Y_15 N_NET15_9 0.00088696f
cc_93 N_Y_3 N_NET15_2 0.00503187f
x_PM_A2O1A1O1Ixp25_ASAP7_75t_R%C VSS C N_MM3_g N_C_1 N_C_4
+ PM_A2O1A1O1Ixp25_ASAP7_75t_R%C
cc_94 N_C_1 N_B_4 0.000906131f
cc_95 N_MM3_g N_MM2_g 0.00330893f
cc_96 N_C_4 N_B_4 0.0053465f
*END of A2O1A1O1Ixp25_ASAP7_75t_R.pxi
.ENDS
*